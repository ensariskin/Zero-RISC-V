`timescale 1ns/1ns

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.09.2025
// Design Name: RV32I Superscalar Processor Core
// Module Name: rv32i_superscalar_core
// Project Name: RV32I Superscalar
// Target Devices: 
// Tool Versions: 
// Description: Top-level module for the RV32I superscalar processor
//              Integrates fetch, buffer, decode, execute, and writeback stages
//              Supports 3-way superscalar execution with out-of-order capabilities
// 
// Dependencies: fetch_buffer_top.sv, multi_fetch.sv, instruction_buffer.sv,
//              decode_stage.sv, execute.sv, mem.sv, write_back.sv
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: 
// - 3-instruction fetch per cycle
// - Variable decode/issue width (1-3 instructions)
// - Branch prediction with fetch optimization
// - Instruction buffer for fetch/decode decoupling
// - Future: Out-of-order execution, register renaming
//////////////////////////////////////////////////////////////////////////////////

module rv32i_superscalar_core #(
    parameter DATA_WIDTH = 32,
    parameter BUFFER_DEPTH = 16,
    parameter REG_FILE_ADDR_WIDTH = 5
)(
    // Clock and Reset
    input  logic clk,
    input  logic reset,
    
    // Instruction Memory Interface (3-port for parallel fetch)
    output logic [DATA_WIDTH-1:0] inst_addr_0, inst_addr_1, inst_addr_2,
    input  logic [DATA_WIDTH-1:0] instruction_i_0, instruction_i_1, instruction_i_2,
    
    // Data Memory Interface (for load/store operations)
    output logic [DATA_WIDTH-1:0] data_addr,
    output logic [DATA_WIDTH-1:0] data_write,
    input  logic [DATA_WIDTH-1:0] data_read,
    output logic data_we,
    output logic [3:0] data_be,
    output logic data_req,
    input  logic data_ack,
    input  logic data_err,
    
    // External Interrupt Interface
    input  logic external_interrupt,
    input  logic timer_interrupt,
    input  logic software_interrupt,
    
    // Debug Interface
    output logic [DATA_WIDTH-1:0] debug_pc,
    output logic [DATA_WIDTH-1:0] debug_instruction,
    output logic debug_valid,
    
    // Performance Counters
    output logic [31:0] perf_cycles,
    output logic [31:0] perf_instructions_fetched,
    output logic [31:0] perf_instructions_executed,
    output logic [31:0] perf_branch_mispredictions,
    output logic [31:0] perf_buffer_stalls,
    
    // Status Outputs
    output logic processor_halted,
    output logic [2:0] current_privilege_mode
);

    localparam D = 1; // Delay for simulation purposes

    // Internal Pipeline Control Signals
    logic pipeline_flush;
    logic pipeline_stall;
    logic decode_bubble;
    
    // Fetch Buffer Interface
    logic [2:0] decode_valid;
    logic [DATA_WIDTH-1:0] fetch_instruction_0, fetch_instruction_1, fetch_instruction_2;
    logic [DATA_WIDTH-1:0] fetch_pc_0, fetch_pc_1, fetch_pc_2;
    logic [DATA_WIDTH-1:0] fetch_imm_0, fetch_imm_1, fetch_imm_2;
    logic fetch_branch_pred_0, fetch_branch_pred_1, fetch_branch_pred_2;
    logic [2:0] decode_ready;
    logic buffer_empty, buffer_full;
    logic [$clog2(BUFFER_DEPTH):0] buffer_occupancy;
    
    // Branch Prediction Interface
    logic [DATA_WIDTH-1:0] bp_pc_0, bp_pc_1, bp_pc_2;
    logic bp_prediction_0, bp_prediction_1, bp_prediction_2;
    logic bp_update_valid_0, bp_update_valid_1, bp_update_valid_2;
    logic [DATA_WIDTH-1:0] bp_update_pc_0, bp_update_pc_1, bp_update_pc_2;
    logic bp_misprediction_0, bp_misprediction_1, bp_misprediction_2;
    logic [DATA_WIDTH-1:0] bp_correct_pc;
    
    // Decode Stage Outputs (3 parallel decode units)
    logic [2:0] decode_valid_out;
    logic [DATA_WIDTH-1:0] decode_data_a_0, decode_data_a_1, decode_data_a_2;
    logic [DATA_WIDTH-1:0] decode_data_b_0, decode_data_b_1, decode_data_b_2;
    logic [DATA_WIDTH-1:0] decode_store_data_0, decode_store_data_1, decode_store_data_2;
    logic [DATA_WIDTH-1:0] decode_pc_0, decode_pc_1, decode_pc_2;
    logic [25:0] decode_control_0, decode_control_1, decode_control_2;
    logic [DATA_WIDTH-1:0] decode_pc_prediction_0, decode_pc_prediction_1, decode_pc_prediction_2;
    logic [2:0] decode_branch_sel_0, decode_branch_sel_1, decode_branch_sel_2;
    logic decode_branch_pred_0, decode_branch_pred_1, decode_branch_pred_2;
    logic [REG_FILE_ADDR_WIDTH-1:0] decode_rs1_0, decode_rs1_1, decode_rs1_2;
    logic [REG_FILE_ADDR_WIDTH-1:0] decode_rs2_0, decode_rs2_1, decode_rs2_2;
    logic [REG_FILE_ADDR_WIDTH-1:0] decode_rd_0, decode_rd_1, decode_rd_2;

    logic [2:0] commit_valid;
    logic [REG_FILE_ADDR_WIDTH-1:0] commit_addr_0;
    logic [REG_FILE_ADDR_WIDTH-1:0] commit_addr_1;
    logic [REG_FILE_ADDR_WIDTH-1:0] commit_addr_2;
    
    // Execute Stage Interface
    logic [2:0] execute_ready;
    logic [2:0] execute_valid_out;
    logic [DATA_WIDTH-1:0] execute_result_0, execute_result_1, execute_result_2;
    logic [REG_FILE_ADDR_WIDTH-1:0] execute_rd_0, execute_rd_1, execute_rd_2;
    logic execute_reg_write_0, execute_reg_write_1, execute_reg_write_2;
    
    // Memory Stage Interface
    logic mem_valid;
    logic [DATA_WIDTH-1:0] mem_result;
    logic [REG_FILE_ADDR_WIDTH-1:0] mem_rd;
    logic mem_reg_write;
    
    // Writeback Stage Interface
    logic [2:0] wb_valid;
    logic [DATA_WIDTH-1:0] wb_data_0, wb_data_1, wb_data_2;
    logic [REG_FILE_ADDR_WIDTH-1:0] wb_rd_0, wb_rd_1, wb_rd_2;
    logic wb_reg_write_0, wb_reg_write_1, wb_reg_write_2;
    
    // Register File Interface (multi-port for superscalar)
    logic [DATA_WIDTH-1:0] rf_read_data_0_0, rf_read_data_0_1; // For instruction 0
    logic [DATA_WIDTH-1:0] rf_read_data_1_0, rf_read_data_1_1; // For instruction 1
    logic [DATA_WIDTH-1:0] rf_read_data_2_0, rf_read_data_2_1; // For instruction 2
    
    // CSR Interface
    logic [11:0] csr_addr;
    logic [DATA_WIDTH-1:0] csr_write_data;
    logic [DATA_WIDTH-1:0] csr_read_data;
    logic csr_write_enable;
    logic csr_read_enable;
    
    // Exception and Interrupt Handling
    logic exception_occurred;
    logic [3:0] exception_cause;
    logic [DATA_WIDTH-1:0] exception_pc;
    logic interrupt_pending;
    
    // Performance Counter Registers
    logic [31:0] cycle_counter;
    logic [31:0] instruction_fetch_counter;
    logic [31:0] instruction_execute_counter;
    logic [31:0] branch_misprediction_counter;
    logic [31:0] buffer_stall_counter;
    
    // Debug and Status Registers
    logic [DATA_WIDTH-1:0] current_pc;
    logic [DATA_WIDTH-1:0] current_instruction;
    logic instruction_valid;
    logic [1:0] privilege_mode;
    logic halted;
    
    //==========================================================================
    // FETCH STAGE (fetch_buffer_top)
    //==========================================================================
    
    fetch_buffer_top #(
        .DATA_WIDTH(DATA_WIDTH),
        .BUFFER_DEPTH(BUFFER_DEPTH)
    ) fetch_buffer_unit (
        .clk(clk),
        .reset(reset),
        
        // Memory interface
        .inst_addr_0(inst_addr_0),
        .instruction_i_0(instruction_i_0),
        .inst_addr_1(inst_addr_1),
        .instruction_i_1(instruction_i_1),
        .inst_addr_2(inst_addr_2),
        .instruction_i_2(instruction_i_2),
        
        // Pipeline control
        .flush(pipeline_flush),
        .buble(pipeline_stall),
        
        // Branch prediction interface
        .pc_value_at_prediction_0(bp_pc_0),
        .branch_prediction_o_0(bp_prediction_0),
        .update_prediction_valid_i_0(bp_update_valid_0),
        .update_prediction_pc_0(bp_update_pc_0),
        .misprediction_0(bp_misprediction_0),
        
        .pc_value_at_prediction_1(bp_pc_1),
        .branch_prediction_o_1(bp_prediction_1),
        .update_prediction_valid_i_1(bp_update_valid_1),
        .update_prediction_pc_1(bp_update_pc_1),
        .misprediction_1(bp_misprediction_1),
        
        .pc_value_at_prediction_2(bp_pc_2),
        .branch_prediction_o_2(bp_prediction_2),
        .update_prediction_valid_i_2(bp_update_valid_2),
        .update_prediction_pc_2(bp_update_pc_2),
        .misprediction_2(bp_misprediction_2),
        
        .correct_pc(bp_correct_pc),
        
        // Output to decode stages
        .decode_valid_o(decode_valid),
        .instruction_o_0(fetch_instruction_0),
        .instruction_o_1(fetch_instruction_1),
        .instruction_o_2(fetch_instruction_2),
        .pc_decode_o_0(fetch_pc_0),
        .pc_decode_o_1(fetch_pc_1),
        .pc_decode_o_2(fetch_pc_2),
        .imm_decode_o_0(fetch_imm_0),
        .imm_decode_o_1(fetch_imm_1),
        .imm_decode_o_2(fetch_imm_2),
        .branch_prediction_decode_o_0(fetch_branch_pred_0),
        .branch_prediction_decode_o_1(fetch_branch_pred_1),
        .branch_prediction_decode_o_2(fetch_branch_pred_2),
        
        // Decode stage ready signals
        .decode_ready_i(decode_ready),
        
        // Status outputs
        .buffer_empty_o(buffer_empty),
        .buffer_full_o(buffer_full),
        .occupancy_o(buffer_occupancy),
        
        // Legacy outputs (not used in superscalar)
        .legacy_instruction_o_0(),
        .legacy_instruction_o_1(),
        .legacy_instruction_o_2(),
        .legacy_imm_o_0(),
        .legacy_imm_o_1(),
        .legacy_imm_o_2(),
        .pc_plus_o()
    );

    
    //==========================================================================
    // ISSUE STAGE (3 parallel decode units with register renaming)
    //==========================================================================
    
    // Create interfaces for issue stage to dispatch stage
    issue_to_dispatch_if #(.DATA_WIDTH(DATA_WIDTH), .PHYS_REG_ADDR_WIDTH(REG_FILE_ADDR_WIDTH+1)) 
        issue_to_dispatch_0_if(), issue_to_dispatch_1_if(), issue_to_dispatch_2_if();
    
    issue_stage #(
        .DATA_WIDTH(DATA_WIDTH),
        .ARCH_REG_ADDR_WIDTH(REG_FILE_ADDR_WIDTH),
        .PHYS_REG_ADDR_WIDTH(REG_FILE_ADDR_WIDTH+1)
    ) issue_stage_unit (
        .clk(clk),
        .reset(reset),
        
        // Pipeline control
        .flush(pipeline_flush),
        .bubble(pipeline_stall),
        
        // Input from fetch/buffer stage
        .decode_valid_i(decode_valid),
        .instruction_i_0(fetch_instruction_0),
        .instruction_i_1(fetch_instruction_1),
        .instruction_i_2(fetch_instruction_2),
        .immediate_i_0(fetch_imm_0),
        .immediate_i_1(fetch_imm_1),
        .immediate_i_2(fetch_imm_2),
        .pc_i_0(fetch_pc_0),
        .pc_i_1(fetch_pc_1),
        .pc_i_2(fetch_pc_2),
        .pc_value_at_prediction_i_0(fetch_pc_0), // Using PC for now
        .pc_value_at_prediction_i_1(fetch_pc_1),
        .pc_value_at_prediction_i_2(fetch_pc_2),
        .branch_prediction_i_0(fetch_branch_pred_0),
        .branch_prediction_i_1(fetch_branch_pred_1),
        .branch_prediction_i_2(fetch_branch_pred_2),
        
        // Ready signal to fetch/buffer stage
        .decode_ready_o(decode_ready),
        
        // ROB commit interface (placeholder for now)
        .commit_addr_0_i(commit_addr_0),
        .commit_addr_1_i(commit_addr_1),
        .commit_addr_2_i(commit_addr_2),
        .commit_valid_i(commit_valid),
        
        // Issue to Dispatch Stage Interfaces
        .issue_to_dispatch_0(issue_to_dispatch_0_if.issue),
        .issue_to_dispatch_1(issue_to_dispatch_1_if.issue),
        .issue_to_dispatch_2(issue_to_dispatch_2_if.issue)
    );
    
    //==========================================================================
    // DISPATCH STAGE (reservation stations + register file)
    //==========================================================================
    
    // Create interfaces for dispatch stage to functional units
    rs_to_exec_if #(.DATA_WIDTH(DATA_WIDTH), .PHYS_REG_ADDR_WIDTH(REG_FILE_ADDR_WIDTH+1)) 
        dispatch_to_alu_0_if(), dispatch_to_alu_1_if(), dispatch_to_alu_2_if();
    
    dispatch_stage #(
        .DATA_WIDTH(DATA_WIDTH),
        .PHYS_REG_ADDR_WIDTH(REG_FILE_ADDR_WIDTH+1),
        .NUM_PHYS_REGS(64)
    ) dispatch_stage_unit (
        .clk(clk),
        .reset(reset),
        
        // Input from Issue Stage
        .issue_to_dispatch_0(issue_to_dispatch_0_if.dispatch),
        .issue_to_dispatch_1(issue_to_dispatch_1_if.dispatch),
        .issue_to_dispatch_2(issue_to_dispatch_2_if.dispatch),
        
        // Output to Functional Units
        .dispatch_to_alu_0(dispatch_to_alu_0_if.reservation_station),
        .dispatch_to_alu_1(dispatch_to_alu_1_if.reservation_station),
        .dispatch_to_alu_2(dispatch_to_alu_2_if.reservation_station),

        .commit_valid(commit_valid),
        .commit_addr_0(commit_addr_0),
        .commit_addr_1(commit_addr_1),
        .commit_addr_2(commit_addr_2)
    );
    
    //==========================================================================
    // EXECUTE STAGE
    //==========================================================================
    
    superscalar_execute_stage #(
        .DATA_WIDTH(DATA_WIDTH)
    ) execute_stage_unit (
        .clk(clk),
        .rst_n(~reset),
        
        // Interface to reservation stations
        .rs_to_exec_0(dispatch_to_alu_0_if.functional_unit),
        .rs_to_exec_1(dispatch_to_alu_1_if.functional_unit),
        .rs_to_exec_2(dispatch_to_alu_2_if.functional_unit)
    );
    
    //==========================================================================
    // TEMPORARY CONNECTIONS (for backward compatibility during transition)
    //==========================================================================
    
    // Extract data from dispatch interfaces for execute stage (temporary)
    assign decode_valid_out[0] = dispatch_to_alu_0_if.issue_valid;
    assign decode_valid_out[1] = dispatch_to_alu_1_if.issue_valid;
    assign decode_valid_out[2] = dispatch_to_alu_2_if.issue_valid;
    
    assign decode_data_a_0 = dispatch_to_alu_0_if.data_a;
    assign decode_data_a_1 = dispatch_to_alu_1_if.data_a;
    assign decode_data_a_2 = dispatch_to_alu_2_if.data_a;
    
    assign decode_data_b_0 = dispatch_to_alu_0_if.data_b;
    assign decode_data_b_1 = dispatch_to_alu_1_if.data_b;
    assign decode_data_b_2 = dispatch_to_alu_2_if.data_b;
    
    assign decode_store_data_0 = dispatch_to_alu_0_if.store_data;  // Now using dedicated store_data signal
    assign decode_store_data_1 = dispatch_to_alu_1_if.store_data;  // Now using dedicated store_data signal
    assign decode_store_data_2 = dispatch_to_alu_2_if.store_data;  // Now using dedicated store_data signal
    
    assign decode_pc_0 = dispatch_to_alu_0_if.pc;                  // Now from rs_to_exec interface
    assign decode_pc_1 = dispatch_to_alu_1_if.pc;                  // Now from rs_to_exec interface
    assign decode_pc_2 = dispatch_to_alu_2_if.pc;                  // Now from rs_to_exec interface
    
    assign decode_control_0 = {15'h0, dispatch_to_alu_0_if.control_signals}; // Now from rs_to_exec interface
    assign decode_control_1 = {15'h0, dispatch_to_alu_1_if.control_signals}; // Now from rs_to_exec interface
    assign decode_control_2 = {15'h0, dispatch_to_alu_2_if.control_signals}; // Now from rs_to_exec interface
    
    assign decode_pc_prediction_0 = dispatch_to_alu_0_if.pc_value_at_prediction;
    assign decode_pc_prediction_1 = dispatch_to_alu_1_if.pc_value_at_prediction;
    assign decode_pc_prediction_2 = dispatch_to_alu_2_if.pc_value_at_prediction;
    
    assign decode_branch_sel_0 = dispatch_to_alu_0_if.branch_sel;
    assign decode_branch_sel_1 = dispatch_to_alu_1_if.branch_sel;
    assign decode_branch_sel_2 = dispatch_to_alu_2_if.branch_sel;
    
    assign decode_branch_pred_0 = dispatch_to_alu_0_if.branch_prediction;
    assign decode_branch_pred_1 = dispatch_to_alu_1_if.branch_prediction;
    assign decode_branch_pred_2 = dispatch_to_alu_2_if.branch_prediction;
    
    // Extract destination registers from rs_to_exec interfaces (convert 6-bit back to 5-bit for now)
    assign decode_rd_0 = dispatch_to_alu_0_if.rd_phys_addr[4:0];
    assign decode_rd_1 = dispatch_to_alu_1_if.rd_phys_addr[4:0];
    assign decode_rd_2 = dispatch_to_alu_2_if.rd_phys_addr[4:0];
    
    //==========================================================================
    // EXECUTE STAGE OUTPUTS (for backward compatibility)
    //==========================================================================
    
    // Extract execute results from interface for temporary compatibility
    assign execute_valid_out = decode_valid_out; // Will be replaced with proper completion signals
    assign execute_result_0 = dispatch_to_alu_0_if.data_result;
    assign execute_result_1 = dispatch_to_alu_1_if.data_result;
    assign execute_result_2 = dispatch_to_alu_2_if.data_result;
    assign execute_rd_0 = decode_rd_0;
    assign execute_rd_1 = decode_rd_1;
    assign execute_rd_2 = decode_rd_2;
    assign execute_reg_write_0 = decode_valid_out[0] & (decode_control_0[0]); // Extract write enable from control
    assign execute_reg_write_1 = decode_valid_out[1] & (decode_control_1[0]); // Extract write enable from control
    assign execute_reg_write_2 = decode_valid_out[2] & (decode_control_2[0]); // Extract write enable from control
    assign execute_ready = 3'b111; // Always ready for now
    
    //==========================================================================
    // MEMORY STAGE (placeholder)
    //==========================================================================
    
    // For now, no memory operations
    // TODO: Implement memory pipeline stage
    assign data_addr = 32'h0;
    assign data_write = 32'h0;
    assign data_we = 1'b0;
    assign data_be = 4'h0;
    assign data_req = 1'b0;
    assign mem_valid = 1'b0;
    assign mem_result = 32'h0;
    assign mem_rd = 5'h0;
    assign mem_reg_write = 1'b0;
    
    //==========================================================================
    // WRITEBACK STAGE (placeholder)
    //==========================================================================
    
    // For now, simple pass-through
    // TODO: Implement proper writeback with register file
    assign wb_valid = execute_valid_out;
    assign wb_data_0 = execute_result_0;
    assign wb_data_1 = execute_result_1;
    assign wb_data_2 = execute_result_2;
    assign wb_rd_0 = execute_rd_0;
    assign wb_rd_1 = execute_rd_1;
    assign wb_rd_2 = execute_rd_2;
    assign wb_reg_write_0 = execute_reg_write_0;
    assign wb_reg_write_1 = execute_reg_write_1;
    assign wb_reg_write_2 = execute_reg_write_2;
    
    //==========================================================================
    // CONTROL AND STATUS
    //==========================================================================
    
    // Pipeline Control Logic
    assign pipeline_flush = 1'b0;
    assign pipeline_stall = 1'b0;
    assign decode_bubble = 1'b0; // Placeholder
    
    // Branch Prediction Updates (placeholder)
    assign bp_update_valid_0 = 1'b0;
    assign bp_update_valid_1 = 1'b0;
    assign bp_update_valid_2 = 1'b0;
    assign bp_update_pc_0 = 32'h0;
    assign bp_update_pc_1 = 32'h0;
    assign bp_update_pc_2 = 32'h0;
    assign bp_misprediction_0 = 1'b0;
    assign bp_misprediction_1 = 1'b0;
    assign bp_misprediction_2 = 1'b0;
    assign bp_correct_pc = 32'h0;
    
    // Exception and Interrupt Handling (placeholder)
    assign exception_occurred = 1'b0;
    assign exception_cause = 4'h0;
    assign exception_pc = 32'h0;
    assign interrupt_pending = external_interrupt | timer_interrupt | software_interrupt;
    
    // CSR Interface (placeholder)
    assign csr_addr = 12'h0;
    assign csr_write_data = 32'h0;
    assign csr_read_data = 32'h0;
    assign csr_write_enable = 1'b0;
    assign csr_read_enable = 1'b0;
    
    //==========================================================================
    // PERFORMANCE COUNTERS
    //==========================================================================
    
    always_ff @(posedge clk or negedge reset) begin
        if (!reset) begin
            cycle_counter <= #D 32'h0;
            instruction_fetch_counter <= #D 32'h0;
            instruction_execute_counter <= #D 32'h0;
            branch_misprediction_counter <= #D 32'h0;
            buffer_stall_counter <= #D 32'h0;
        end else begin
            cycle_counter <= #D cycle_counter + 1;
            
            // Count fetched instructions
            instruction_fetch_counter <= #D instruction_fetch_counter + 
                                       decode_valid[0] + decode_valid[1] + decode_valid[2];
            
            // Count executed instructions
            instruction_execute_counter <= #D instruction_execute_counter + 
                                         execute_valid_out[0] + execute_valid_out[1] + execute_valid_out[2];
            
            // Count branch mispredictions
            if (bp_misprediction_0 | bp_misprediction_1 | bp_misprediction_2) begin
                branch_misprediction_counter <= #D branch_misprediction_counter + 1;
            end
            
            // Count buffer stalls
            if (buffer_full) begin
                buffer_stall_counter <= #D buffer_stall_counter + 1;
            end
        end
    end
    
    //==========================================================================
    // DEBUG AND STATUS OUTPUTS
    //==========================================================================
    
    // Debug interface
    assign debug_pc = inst_addr_0;
    assign debug_instruction = fetch_instruction_0;
    assign debug_valid = decode_valid[0];
    
    // Status outputs
    assign processor_halted = halted;
    assign current_privilege_mode = {1'b0, privilege_mode};
    
    // Performance counter outputs
    assign perf_cycles = cycle_counter;
    assign perf_instructions_fetched = instruction_fetch_counter;
    assign perf_instructions_executed = instruction_execute_counter;
    assign perf_branch_mispredictions = branch_misprediction_counter;
    assign perf_buffer_stalls = buffer_stall_counter;
    
    // Status registers
    assign halted = 1'b0; // Placeholder
    assign privilege_mode = 2'b11; // Machine mode
    assign current_pc = fetch_pc_0;
    assign current_instruction = fetch_instruction_0;
    assign instruction_valid = decode_valid[0];

endmodule
