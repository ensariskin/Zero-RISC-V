// Final fault injection target list (deduplicated & cleaned)
// Signals under 'dv_top.dut.', excluding clk/reset/tracer, compacted by bit-range

//parameter int NUM_FAULT_TARGETS = 1652;
logic [31:0] fi_targets[1652];

// Target aliases
alias fi_targets[0] = dv_top.dut.DF.A_sel;
alias fi_targets[1] = dv_top.dut.DF.B_sel;
alias fi_targets[2] = dv_top.dut.DF.MB;
alias fi_targets[3] = dv_top.dut.DF.RA;
alias fi_targets[4] = dv_top.dut.DF.RA_RD_MEM;
alias fi_targets[5] = dv_top.dut.DF.RA_RD_MEM_exor;
alias fi_targets[6] = dv_top.dut.DF.RA_RD_WB;
alias fi_targets[7] = dv_top.dut.DF.RA_RD_WB_exor;
alias fi_targets[8] = dv_top.dut.DF.RB;
alias fi_targets[9] = dv_top.dut.DF.RB_RD_MEM;
alias fi_targets[10] = dv_top.dut.DF.RB_RD_MEM_exor;
alias fi_targets[11] = dv_top.dut.DF.RB_RD_WB;
alias fi_targets[12] = dv_top.dut.DF.RB_RD_WB_exor;
alias fi_targets[13] = dv_top.dut.DF.RD_MEM;
alias fi_targets[14] = dv_top.dut.DF.RD_WB;
alias fi_targets[15] = dv_top.dut.DF.WE_MEM;
alias fi_targets[16] = dv_top.dut.DF.WE_WB;
alias fi_targets[17] = dv_top.dut.DF.store_data_sel;
alias fi_targets[18] = dv_top.dut.EX.branch_controller.MUX.addr;
alias fi_targets[19] = dv_top.dut.EX.branch_controller.MUX.data_in;
alias fi_targets[20] = dv_top.dut.EX.branch_controller.MUX.data_out;
alias fi_targets[21] = dv_top.dut.EX.branch_controller.MUX.inner_data;
alias fi_targets[22] = dv_top.dut.EX.branch_controller.Branch_sel;
alias fi_targets[23] = dv_top.dut.EX.branch_controller.JALR;
alias fi_targets[24] = dv_top.dut.EX.branch_controller.MPC;
alias fi_targets[25] = dv_top.dut.EX.branch_controller.N;
alias fi_targets[26] = dv_top.dut.EX.branch_controller.Z;
alias fi_targets[27] = dv_top.dut.EX.dat_b_mux.addr;
alias fi_targets[28] = dv_top.dut.EX.dat_b_mux.data_in;
alias fi_targets[29] = dv_top.dut.EX.dat_b_mux.data_out;
alias fi_targets[30] = dv_top.dut.EX.dat_b_mux.inner_data;
alias fi_targets[31] = dv_top.dut.EX.data_a_mux.addr;
alias fi_targets[32] = dv_top.dut.EX.data_a_mux.data_in;
alias fi_targets[33] = dv_top.dut.EX.data_a_mux.data_out;
alias fi_targets[34] = dv_top.dut.EX.data_a_mux.inner_data;
alias fi_targets[35] = dv_top.dut.EX.data_store_mux.addr;
alias fi_targets[36] = dv_top.dut.EX.data_store_mux.data_in;
alias fi_targets[37] = dv_top.dut.EX.data_store_mux.data_out;
alias fi_targets[38] = dv_top.dut.EX.data_store_mux.inner_data;
alias fi_targets[39] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.half_adder_1.cout;
alias fi_targets[40] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.half_adder_1.s;
alias fi_targets[41] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.half_adder_1.x;
alias fi_targets[42] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.half_adder_1.y;
alias fi_targets[43] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.half_adder_2.cout;
alias fi_targets[44] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.half_adder_2.s;
alias fi_targets[45] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.half_adder_2.x;
alias fi_targets[46] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.half_adder_2.y;
alias fi_targets[47] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.c0;
alias fi_targets[48] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.c1;
alias fi_targets[49] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.ci;
alias fi_targets[50] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.cout;
alias fi_targets[51] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.s;
alias fi_targets[52] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.s0;
alias fi_targets[53] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.x;
alias fi_targets[54] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[0].full_adder.y;
alias fi_targets[55] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.half_adder_1.cout;
alias fi_targets[56] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.half_adder_1.s;
alias fi_targets[57] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.half_adder_1.x;
alias fi_targets[58] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.half_adder_1.y;
alias fi_targets[59] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.half_adder_2.cout;
alias fi_targets[60] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.half_adder_2.s;
alias fi_targets[61] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.half_adder_2.x;
alias fi_targets[62] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.half_adder_2.y;
alias fi_targets[63] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.c0;
alias fi_targets[64] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.c1;
alias fi_targets[65] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.ci;
alias fi_targets[66] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.cout;
alias fi_targets[67] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.s;
alias fi_targets[68] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.s0;
alias fi_targets[69] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.x;
alias fi_targets[70] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[10].full_adder.y;
alias fi_targets[71] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.half_adder_1.cout;
alias fi_targets[72] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.half_adder_1.s;
alias fi_targets[73] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.half_adder_1.x;
alias fi_targets[74] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.half_adder_1.y;
alias fi_targets[75] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.half_adder_2.cout;
alias fi_targets[76] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.half_adder_2.s;
alias fi_targets[77] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.half_adder_2.x;
alias fi_targets[78] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.half_adder_2.y;
alias fi_targets[79] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.c0;
alias fi_targets[80] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.c1;
alias fi_targets[81] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.ci;
alias fi_targets[82] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.cout;
alias fi_targets[83] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.s;
alias fi_targets[84] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.s0;
alias fi_targets[85] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.x;
alias fi_targets[86] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[11].full_adder.y;
alias fi_targets[87] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.half_adder_1.cout;
alias fi_targets[88] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.half_adder_1.s;
alias fi_targets[89] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.half_adder_1.x;
alias fi_targets[90] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.half_adder_1.y;
alias fi_targets[91] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.half_adder_2.cout;
alias fi_targets[92] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.half_adder_2.s;
alias fi_targets[93] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.half_adder_2.x;
alias fi_targets[94] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.half_adder_2.y;
alias fi_targets[95] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.c0;
alias fi_targets[96] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.c1;
alias fi_targets[97] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.ci;
alias fi_targets[98] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.cout;
alias fi_targets[99] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.s;
alias fi_targets[100] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.s0;
alias fi_targets[101] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.x;
alias fi_targets[102] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[12].full_adder.y;
alias fi_targets[103] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.half_adder_1.cout;
alias fi_targets[104] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.half_adder_1.s;
alias fi_targets[105] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.half_adder_1.x;
alias fi_targets[106] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.half_adder_1.y;
alias fi_targets[107] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.half_adder_2.cout;
alias fi_targets[108] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.half_adder_2.s;
alias fi_targets[109] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.half_adder_2.x;
alias fi_targets[110] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.half_adder_2.y;
alias fi_targets[111] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.c0;
alias fi_targets[112] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.c1;
alias fi_targets[113] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.ci;
alias fi_targets[114] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.cout;
alias fi_targets[115] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.s;
alias fi_targets[116] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.s0;
alias fi_targets[117] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.x;
alias fi_targets[118] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[13].full_adder.y;
alias fi_targets[119] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.half_adder_1.cout;
alias fi_targets[120] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.half_adder_1.s;
alias fi_targets[121] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.half_adder_1.x;
alias fi_targets[122] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.half_adder_1.y;
alias fi_targets[123] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.half_adder_2.cout;
alias fi_targets[124] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.half_adder_2.s;
alias fi_targets[125] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.half_adder_2.x;
alias fi_targets[126] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.half_adder_2.y;
alias fi_targets[127] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.c0;
alias fi_targets[128] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.c1;
alias fi_targets[129] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.ci;
alias fi_targets[130] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.cout;
alias fi_targets[131] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.s;
alias fi_targets[132] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.s0;
alias fi_targets[133] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.x;
alias fi_targets[134] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[14].full_adder.y;
alias fi_targets[135] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.half_adder_1.cout;
alias fi_targets[136] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.half_adder_1.s;
alias fi_targets[137] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.half_adder_1.x;
alias fi_targets[138] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.half_adder_1.y;
alias fi_targets[139] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.half_adder_2.cout;
alias fi_targets[140] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.half_adder_2.s;
alias fi_targets[141] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.half_adder_2.x;
alias fi_targets[142] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.half_adder_2.y;
alias fi_targets[143] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.c0;
alias fi_targets[144] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.c1;
alias fi_targets[145] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.ci;
alias fi_targets[146] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.cout;
alias fi_targets[147] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.s;
alias fi_targets[148] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.s0;
alias fi_targets[149] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.x;
alias fi_targets[150] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[15].full_adder.y;
alias fi_targets[151] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.half_adder_1.cout;
alias fi_targets[152] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.half_adder_1.s;
alias fi_targets[153] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.half_adder_1.x;
alias fi_targets[154] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.half_adder_1.y;
alias fi_targets[155] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.half_adder_2.cout;
alias fi_targets[156] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.half_adder_2.s;
alias fi_targets[157] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.half_adder_2.x;
alias fi_targets[158] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.half_adder_2.y;
alias fi_targets[159] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.c0;
alias fi_targets[160] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.c1;
alias fi_targets[161] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.ci;
alias fi_targets[162] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.cout;
alias fi_targets[163] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.s;
alias fi_targets[164] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.s0;
alias fi_targets[165] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.x;
alias fi_targets[166] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[16].full_adder.y;
alias fi_targets[167] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.half_adder_1.cout;
alias fi_targets[168] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.half_adder_1.s;
alias fi_targets[169] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.half_adder_1.x;
alias fi_targets[170] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.half_adder_1.y;
alias fi_targets[171] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.half_adder_2.cout;
alias fi_targets[172] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.half_adder_2.s;
alias fi_targets[173] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.half_adder_2.x;
alias fi_targets[174] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.half_adder_2.y;
alias fi_targets[175] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.c0;
alias fi_targets[176] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.c1;
alias fi_targets[177] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.ci;
alias fi_targets[178] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.cout;
alias fi_targets[179] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.s;
alias fi_targets[180] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.s0;
alias fi_targets[181] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.x;
alias fi_targets[182] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[17].full_adder.y;
alias fi_targets[183] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.half_adder_1.cout;
alias fi_targets[184] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.half_adder_1.s;
alias fi_targets[185] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.half_adder_1.x;
alias fi_targets[186] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.half_adder_1.y;
alias fi_targets[187] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.half_adder_2.cout;
alias fi_targets[188] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.half_adder_2.s;
alias fi_targets[189] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.half_adder_2.x;
alias fi_targets[190] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.half_adder_2.y;
alias fi_targets[191] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.c0;
alias fi_targets[192] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.c1;
alias fi_targets[193] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.ci;
alias fi_targets[194] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.cout;
alias fi_targets[195] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.s;
alias fi_targets[196] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.s0;
alias fi_targets[197] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.x;
alias fi_targets[198] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[18].full_adder.y;
alias fi_targets[199] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.half_adder_1.cout;
alias fi_targets[200] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.half_adder_1.s;
alias fi_targets[201] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.half_adder_1.x;
alias fi_targets[202] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.half_adder_1.y;
alias fi_targets[203] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.half_adder_2.cout;
alias fi_targets[204] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.half_adder_2.s;
alias fi_targets[205] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.half_adder_2.x;
alias fi_targets[206] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.half_adder_2.y;
alias fi_targets[207] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.c0;
alias fi_targets[208] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.c1;
alias fi_targets[209] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.ci;
alias fi_targets[210] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.cout;
alias fi_targets[211] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.s;
alias fi_targets[212] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.s0;
alias fi_targets[213] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.x;
alias fi_targets[214] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[19].full_adder.y;
alias fi_targets[215] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.half_adder_1.cout;
alias fi_targets[216] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.half_adder_1.s;
alias fi_targets[217] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.half_adder_1.x;
alias fi_targets[218] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.half_adder_1.y;
alias fi_targets[219] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.half_adder_2.cout;
alias fi_targets[220] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.half_adder_2.s;
alias fi_targets[221] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.half_adder_2.x;
alias fi_targets[222] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.half_adder_2.y;
alias fi_targets[223] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.c0;
alias fi_targets[224] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.c1;
alias fi_targets[225] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.ci;
alias fi_targets[226] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.cout;
alias fi_targets[227] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.s;
alias fi_targets[228] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.s0;
alias fi_targets[229] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.x;
alias fi_targets[230] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[1].full_adder.y;
alias fi_targets[231] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.half_adder_1.cout;
alias fi_targets[232] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.half_adder_1.s;
alias fi_targets[233] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.half_adder_1.x;
alias fi_targets[234] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.half_adder_1.y;
alias fi_targets[235] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.half_adder_2.cout;
alias fi_targets[236] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.half_adder_2.s;
alias fi_targets[237] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.half_adder_2.x;
alias fi_targets[238] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.half_adder_2.y;
alias fi_targets[239] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.c0;
alias fi_targets[240] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.c1;
alias fi_targets[241] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.ci;
alias fi_targets[242] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.cout;
alias fi_targets[243] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.s;
alias fi_targets[244] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.s0;
alias fi_targets[245] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.x;
alias fi_targets[246] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[20].full_adder.y;
alias fi_targets[247] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.half_adder_1.cout;
alias fi_targets[248] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.half_adder_1.s;
alias fi_targets[249] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.half_adder_1.x;
alias fi_targets[250] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.half_adder_1.y;
alias fi_targets[251] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.half_adder_2.cout;
alias fi_targets[252] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.half_adder_2.s;
alias fi_targets[253] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.half_adder_2.x;
alias fi_targets[254] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.half_adder_2.y;
alias fi_targets[255] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.c0;
alias fi_targets[256] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.c1;
alias fi_targets[257] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.ci;
alias fi_targets[258] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.cout;
alias fi_targets[259] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.s;
alias fi_targets[260] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.s0;
alias fi_targets[261] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.x;
alias fi_targets[262] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[21].full_adder.y;
alias fi_targets[263] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.half_adder_1.cout;
alias fi_targets[264] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.half_adder_1.s;
alias fi_targets[265] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.half_adder_1.x;
alias fi_targets[266] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.half_adder_1.y;
alias fi_targets[267] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.half_adder_2.cout;
alias fi_targets[268] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.half_adder_2.s;
alias fi_targets[269] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.half_adder_2.x;
alias fi_targets[270] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.half_adder_2.y;
alias fi_targets[271] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.c0;
alias fi_targets[272] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.c1;
alias fi_targets[273] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.ci;
alias fi_targets[274] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.cout;
alias fi_targets[275] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.s;
alias fi_targets[276] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.s0;
alias fi_targets[277] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.x;
alias fi_targets[278] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[22].full_adder.y;
alias fi_targets[279] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.half_adder_1.cout;
alias fi_targets[280] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.half_adder_1.s;
alias fi_targets[281] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.half_adder_1.x;
alias fi_targets[282] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.half_adder_1.y;
alias fi_targets[283] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.half_adder_2.cout;
alias fi_targets[284] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.half_adder_2.s;
alias fi_targets[285] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.half_adder_2.x;
alias fi_targets[286] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.half_adder_2.y;
alias fi_targets[287] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.c0;
alias fi_targets[288] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.c1;
alias fi_targets[289] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.ci;
alias fi_targets[290] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.cout;
alias fi_targets[291] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.s;
alias fi_targets[292] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.s0;
alias fi_targets[293] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.x;
alias fi_targets[294] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[23].full_adder.y;
alias fi_targets[295] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.half_adder_1.cout;
alias fi_targets[296] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.half_adder_1.s;
alias fi_targets[297] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.half_adder_1.x;
alias fi_targets[298] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.half_adder_1.y;
alias fi_targets[299] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.half_adder_2.cout;
alias fi_targets[300] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.half_adder_2.s;
alias fi_targets[301] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.half_adder_2.x;
alias fi_targets[302] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.half_adder_2.y;
alias fi_targets[303] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.c0;
alias fi_targets[304] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.c1;
alias fi_targets[305] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.ci;
alias fi_targets[306] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.cout;
alias fi_targets[307] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.s;
alias fi_targets[308] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.s0;
alias fi_targets[309] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.x;
alias fi_targets[310] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[24].full_adder.y;
alias fi_targets[311] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.half_adder_1.cout;
alias fi_targets[312] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.half_adder_1.s;
alias fi_targets[313] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.half_adder_1.x;
alias fi_targets[314] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.half_adder_1.y;
alias fi_targets[315] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.half_adder_2.cout;
alias fi_targets[316] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.half_adder_2.s;
alias fi_targets[317] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.half_adder_2.x;
alias fi_targets[318] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.half_adder_2.y;
alias fi_targets[319] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.c0;
alias fi_targets[320] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.c1;
alias fi_targets[321] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.ci;
alias fi_targets[322] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.cout;
alias fi_targets[323] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.s;
alias fi_targets[324] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.s0;
alias fi_targets[325] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.x;
alias fi_targets[326] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[25].full_adder.y;
alias fi_targets[327] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.half_adder_1.cout;
alias fi_targets[328] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.half_adder_1.s;
alias fi_targets[329] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.half_adder_1.x;
alias fi_targets[330] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.half_adder_1.y;
alias fi_targets[331] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.half_adder_2.cout;
alias fi_targets[332] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.half_adder_2.s;
alias fi_targets[333] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.half_adder_2.x;
alias fi_targets[334] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.half_adder_2.y;
alias fi_targets[335] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.c0;
alias fi_targets[336] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.c1;
alias fi_targets[337] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.ci;
alias fi_targets[338] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.cout;
alias fi_targets[339] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.s;
alias fi_targets[340] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.s0;
alias fi_targets[341] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.x;
alias fi_targets[342] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[26].full_adder.y;
alias fi_targets[343] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.half_adder_1.cout;
alias fi_targets[344] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.half_adder_1.s;
alias fi_targets[345] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.half_adder_1.x;
alias fi_targets[346] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.half_adder_1.y;
alias fi_targets[347] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.half_adder_2.cout;
alias fi_targets[348] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.half_adder_2.s;
alias fi_targets[349] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.half_adder_2.x;
alias fi_targets[350] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.half_adder_2.y;
alias fi_targets[351] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.c0;
alias fi_targets[352] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.c1;
alias fi_targets[353] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.ci;
alias fi_targets[354] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.cout;
alias fi_targets[355] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.s;
alias fi_targets[356] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.s0;
alias fi_targets[357] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.x;
alias fi_targets[358] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[27].full_adder.y;
alias fi_targets[359] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.half_adder_1.cout;
alias fi_targets[360] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.half_adder_1.s;
alias fi_targets[361] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.half_adder_1.x;
alias fi_targets[362] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.half_adder_1.y;
alias fi_targets[363] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.half_adder_2.cout;
alias fi_targets[364] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.half_adder_2.s;
alias fi_targets[365] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.half_adder_2.x;
alias fi_targets[366] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.half_adder_2.y;
alias fi_targets[367] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.c0;
alias fi_targets[368] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.c1;
alias fi_targets[369] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.ci;
alias fi_targets[370] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.cout;
alias fi_targets[371] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.s;
alias fi_targets[372] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.s0;
alias fi_targets[373] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.x;
alias fi_targets[374] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[28].full_adder.y;
alias fi_targets[375] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.half_adder_1.cout;
alias fi_targets[376] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.half_adder_1.s;
alias fi_targets[377] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.half_adder_1.x;
alias fi_targets[378] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.half_adder_1.y;
alias fi_targets[379] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.half_adder_2.cout;
alias fi_targets[380] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.half_adder_2.s;
alias fi_targets[381] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.half_adder_2.x;
alias fi_targets[382] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.half_adder_2.y;
alias fi_targets[383] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.c0;
alias fi_targets[384] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.c1;
alias fi_targets[385] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.ci;
alias fi_targets[386] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.cout;
alias fi_targets[387] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.s;
alias fi_targets[388] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.s0;
alias fi_targets[389] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.x;
alias fi_targets[390] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[29].full_adder.y;
alias fi_targets[391] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.half_adder_1.cout;
alias fi_targets[392] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.half_adder_1.s;
alias fi_targets[393] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.half_adder_1.x;
alias fi_targets[394] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.half_adder_1.y;
alias fi_targets[395] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.half_adder_2.cout;
alias fi_targets[396] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.half_adder_2.s;
alias fi_targets[397] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.half_adder_2.x;
alias fi_targets[398] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.half_adder_2.y;
alias fi_targets[399] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.c0;
alias fi_targets[400] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.c1;
alias fi_targets[401] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.ci;
alias fi_targets[402] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.cout;
alias fi_targets[403] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.s;
alias fi_targets[404] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.s0;
alias fi_targets[405] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.x;
alias fi_targets[406] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[2].full_adder.y;
alias fi_targets[407] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.half_adder_1.cout;
alias fi_targets[408] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.half_adder_1.s;
alias fi_targets[409] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.half_adder_1.x;
alias fi_targets[410] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.half_adder_1.y;
alias fi_targets[411] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.half_adder_2.cout;
alias fi_targets[412] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.half_adder_2.s;
alias fi_targets[413] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.half_adder_2.x;
alias fi_targets[414] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.half_adder_2.y;
alias fi_targets[415] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.c0;
alias fi_targets[416] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.c1;
alias fi_targets[417] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.ci;
alias fi_targets[418] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.cout;
alias fi_targets[419] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.s;
alias fi_targets[420] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.s0;
alias fi_targets[421] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.x;
alias fi_targets[422] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[30].full_adder.y;
alias fi_targets[423] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.half_adder_1.cout;
alias fi_targets[424] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.half_adder_1.s;
alias fi_targets[425] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.half_adder_1.x;
alias fi_targets[426] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.half_adder_1.y;
alias fi_targets[427] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.half_adder_2.cout;
alias fi_targets[428] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.half_adder_2.s;
alias fi_targets[429] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.half_adder_2.x;
alias fi_targets[430] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.half_adder_2.y;
alias fi_targets[431] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.c0;
alias fi_targets[432] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.c1;
alias fi_targets[433] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.ci;
alias fi_targets[434] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.cout;
alias fi_targets[435] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.s;
alias fi_targets[436] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.s0;
alias fi_targets[437] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.x;
alias fi_targets[438] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[31].full_adder.y;
alias fi_targets[439] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.half_adder_1.cout;
alias fi_targets[440] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.half_adder_1.s;
alias fi_targets[441] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.half_adder_1.x;
alias fi_targets[442] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.half_adder_1.y;
alias fi_targets[443] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.half_adder_2.cout;
alias fi_targets[444] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.half_adder_2.s;
alias fi_targets[445] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.half_adder_2.x;
alias fi_targets[446] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.half_adder_2.y;
alias fi_targets[447] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.c0;
alias fi_targets[448] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.c1;
alias fi_targets[449] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.ci;
alias fi_targets[450] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.cout;
alias fi_targets[451] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.s;
alias fi_targets[452] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.s0;
alias fi_targets[453] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.x;
alias fi_targets[454] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[3].full_adder.y;
alias fi_targets[455] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.half_adder_1.cout;
alias fi_targets[456] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.half_adder_1.s;
alias fi_targets[457] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.half_adder_1.x;
alias fi_targets[458] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.half_adder_1.y;
alias fi_targets[459] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.half_adder_2.cout;
alias fi_targets[460] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.half_adder_2.s;
alias fi_targets[461] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.half_adder_2.x;
alias fi_targets[462] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.half_adder_2.y;
alias fi_targets[463] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.c0;
alias fi_targets[464] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.c1;
alias fi_targets[465] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.ci;
alias fi_targets[466] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.cout;
alias fi_targets[467] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.s;
alias fi_targets[468] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.s0;
alias fi_targets[469] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.x;
alias fi_targets[470] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[4].full_adder.y;
alias fi_targets[471] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.half_adder_1.cout;
alias fi_targets[472] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.half_adder_1.s;
alias fi_targets[473] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.half_adder_1.x;
alias fi_targets[474] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.half_adder_1.y;
alias fi_targets[475] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.half_adder_2.cout;
alias fi_targets[476] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.half_adder_2.s;
alias fi_targets[477] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.half_adder_2.x;
alias fi_targets[478] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.half_adder_2.y;
alias fi_targets[479] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.c0;
alias fi_targets[480] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.c1;
alias fi_targets[481] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.ci;
alias fi_targets[482] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.cout;
alias fi_targets[483] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.s;
alias fi_targets[484] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.s0;
alias fi_targets[485] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.x;
alias fi_targets[486] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[5].full_adder.y;
alias fi_targets[487] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.half_adder_1.cout;
alias fi_targets[488] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.half_adder_1.s;
alias fi_targets[489] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.half_adder_1.x;
alias fi_targets[490] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.half_adder_1.y;
alias fi_targets[491] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.half_adder_2.cout;
alias fi_targets[492] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.half_adder_2.s;
alias fi_targets[493] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.half_adder_2.x;
alias fi_targets[494] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.half_adder_2.y;
alias fi_targets[495] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.c0;
alias fi_targets[496] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.c1;
alias fi_targets[497] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.ci;
alias fi_targets[498] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.cout;
alias fi_targets[499] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.s;
alias fi_targets[500] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.s0;
alias fi_targets[501] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.x;
alias fi_targets[502] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[6].full_adder.y;
alias fi_targets[503] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.half_adder_1.cout;
alias fi_targets[504] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.half_adder_1.s;
alias fi_targets[505] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.half_adder_1.x;
alias fi_targets[506] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.half_adder_1.y;
alias fi_targets[507] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.half_adder_2.cout;
alias fi_targets[508] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.half_adder_2.s;
alias fi_targets[509] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.half_adder_2.x;
alias fi_targets[510] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.half_adder_2.y;
alias fi_targets[511] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.c0;
alias fi_targets[512] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.c1;
alias fi_targets[513] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.ci;
alias fi_targets[514] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.cout;
alias fi_targets[515] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.s;
alias fi_targets[516] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.s0;
alias fi_targets[517] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.x;
alias fi_targets[518] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[7].full_adder.y;
alias fi_targets[519] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.half_adder_1.cout;
alias fi_targets[520] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.half_adder_1.s;
alias fi_targets[521] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.half_adder_1.x;
alias fi_targets[522] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.half_adder_1.y;
alias fi_targets[523] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.half_adder_2.cout;
alias fi_targets[524] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.half_adder_2.s;
alias fi_targets[525] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.half_adder_2.x;
alias fi_targets[526] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.half_adder_2.y;
alias fi_targets[527] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.c0;
alias fi_targets[528] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.c1;
alias fi_targets[529] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.ci;
alias fi_targets[530] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.cout;
alias fi_targets[531] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.s;
alias fi_targets[532] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.s0;
alias fi_targets[533] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.x;
alias fi_targets[534] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[8].full_adder.y;
alias fi_targets[535] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.half_adder_1.cout;
alias fi_targets[536] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.half_adder_1.s;
alias fi_targets[537] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.half_adder_1.x;
alias fi_targets[538] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.half_adder_1.y;
alias fi_targets[539] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.half_adder_2.cout;
alias fi_targets[540] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.half_adder_2.s;
alias fi_targets[541] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.half_adder_2.x;
alias fi_targets[542] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.half_adder_2.y;
alias fi_targets[543] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.c0;
alias fi_targets[544] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.c1;
alias fi_targets[545] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.ci;
alias fi_targets[546] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.cout;
alias fi_targets[547] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.s;
alias fi_targets[548] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.s0;
alias fi_targets[549] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.x;
alias fi_targets[550] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.genblk1[9].full_adder.y;
alias fi_targets[551] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.c;
alias fi_targets[552] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.ci;
alias fi_targets[553] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.cout;
alias fi_targets[554] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.s;
alias fi_targets[555] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.x;
alias fi_targets[556] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.final_stage.y;
alias fi_targets[557] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.half_adder_1.cout;
alias fi_targets[558] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.half_adder_1.s;
alias fi_targets[559] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.half_adder_1.x;
alias fi_targets[560] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.half_adder_1.y;
alias fi_targets[561] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.half_adder_2.cout;
alias fi_targets[562] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.half_adder_2.s;
alias fi_targets[563] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.half_adder_2.x;
alias fi_targets[564] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.half_adder_2.y;
alias fi_targets[565] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.c0;
alias fi_targets[566] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.c1;
alias fi_targets[567] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.ci;
alias fi_targets[568] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.cout;
alias fi_targets[569] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.s;
alias fi_targets[570] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.s0;
alias fi_targets[571] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.x;
alias fi_targets[572] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[0].first_stage.y;
alias fi_targets[573] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.half_adder_1.cout;
alias fi_targets[574] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.half_adder_1.s;
alias fi_targets[575] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.half_adder_1.x;
alias fi_targets[576] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.half_adder_1.y;
alias fi_targets[577] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.half_adder_2.cout;
alias fi_targets[578] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.half_adder_2.s;
alias fi_targets[579] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.half_adder_2.x;
alias fi_targets[580] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.half_adder_2.y;
alias fi_targets[581] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.c0;
alias fi_targets[582] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.c1;
alias fi_targets[583] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.ci;
alias fi_targets[584] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.cout;
alias fi_targets[585] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.s;
alias fi_targets[586] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.s0;
alias fi_targets[587] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.x;
alias fi_targets[588] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[10].first_stage.y;
alias fi_targets[589] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.half_adder_1.cout;
alias fi_targets[590] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.half_adder_1.s;
alias fi_targets[591] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.half_adder_1.x;
alias fi_targets[592] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.half_adder_1.y;
alias fi_targets[593] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.half_adder_2.cout;
alias fi_targets[594] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.half_adder_2.s;
alias fi_targets[595] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.half_adder_2.x;
alias fi_targets[596] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.half_adder_2.y;
alias fi_targets[597] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.c0;
alias fi_targets[598] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.c1;
alias fi_targets[599] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.ci;
alias fi_targets[600] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.cout;
alias fi_targets[601] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.s;
alias fi_targets[602] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.s0;
alias fi_targets[603] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.x;
alias fi_targets[604] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[11].first_stage.y;
alias fi_targets[605] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.half_adder_1.cout;
alias fi_targets[606] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.half_adder_1.s;
alias fi_targets[607] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.half_adder_1.x;
alias fi_targets[608] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.half_adder_1.y;
alias fi_targets[609] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.half_adder_2.cout;
alias fi_targets[610] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.half_adder_2.s;
alias fi_targets[611] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.half_adder_2.x;
alias fi_targets[612] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.half_adder_2.y;
alias fi_targets[613] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.c0;
alias fi_targets[614] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.c1;
alias fi_targets[615] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.ci;
alias fi_targets[616] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.cout;
alias fi_targets[617] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.s;
alias fi_targets[618] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.s0;
alias fi_targets[619] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.x;
alias fi_targets[620] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[12].first_stage.y;
alias fi_targets[621] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.half_adder_1.cout;
alias fi_targets[622] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.half_adder_1.s;
alias fi_targets[623] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.half_adder_1.x;
alias fi_targets[624] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.half_adder_1.y;
alias fi_targets[625] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.half_adder_2.cout;
alias fi_targets[626] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.half_adder_2.s;
alias fi_targets[627] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.half_adder_2.x;
alias fi_targets[628] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.half_adder_2.y;
alias fi_targets[629] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.c0;
alias fi_targets[630] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.c1;
alias fi_targets[631] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.ci;
alias fi_targets[632] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.cout;
alias fi_targets[633] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.s;
alias fi_targets[634] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.s0;
alias fi_targets[635] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.x;
alias fi_targets[636] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[13].first_stage.y;
alias fi_targets[637] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.half_adder_1.cout;
alias fi_targets[638] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.half_adder_1.s;
alias fi_targets[639] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.half_adder_1.x;
alias fi_targets[640] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.half_adder_1.y;
alias fi_targets[641] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.half_adder_2.cout;
alias fi_targets[642] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.half_adder_2.s;
alias fi_targets[643] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.half_adder_2.x;
alias fi_targets[644] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.half_adder_2.y;
alias fi_targets[645] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.c0;
alias fi_targets[646] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.c1;
alias fi_targets[647] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.ci;
alias fi_targets[648] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.cout;
alias fi_targets[649] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.s;
alias fi_targets[650] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.s0;
alias fi_targets[651] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.x;
alias fi_targets[652] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[14].first_stage.y;
alias fi_targets[653] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.half_adder_1.cout;
alias fi_targets[654] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.half_adder_1.s;
alias fi_targets[655] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.half_adder_1.x;
alias fi_targets[656] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.half_adder_1.y;
alias fi_targets[657] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.half_adder_2.cout;
alias fi_targets[658] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.half_adder_2.s;
alias fi_targets[659] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.half_adder_2.x;
alias fi_targets[660] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.half_adder_2.y;
alias fi_targets[661] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.c0;
alias fi_targets[662] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.c1;
alias fi_targets[663] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.ci;
alias fi_targets[664] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.cout;
alias fi_targets[665] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.s;
alias fi_targets[666] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.s0;
alias fi_targets[667] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.x;
alias fi_targets[668] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[15].first_stage.y;
alias fi_targets[669] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.half_adder_1.cout;
alias fi_targets[670] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.half_adder_1.s;
alias fi_targets[671] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.half_adder_1.x;
alias fi_targets[672] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.half_adder_1.y;
alias fi_targets[673] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.half_adder_2.cout;
alias fi_targets[674] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.half_adder_2.s;
alias fi_targets[675] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.half_adder_2.x;
alias fi_targets[676] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.half_adder_2.y;
alias fi_targets[677] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.c0;
alias fi_targets[678] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.c1;
alias fi_targets[679] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.ci;
alias fi_targets[680] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.cout;
alias fi_targets[681] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.s;
alias fi_targets[682] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.s0;
alias fi_targets[683] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.x;
alias fi_targets[684] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[16].first_stage.y;
alias fi_targets[685] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.half_adder_1.cout;
alias fi_targets[686] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.half_adder_1.s;
alias fi_targets[687] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.half_adder_1.x;
alias fi_targets[688] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.half_adder_1.y;
alias fi_targets[689] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.half_adder_2.cout;
alias fi_targets[690] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.half_adder_2.s;
alias fi_targets[691] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.half_adder_2.x;
alias fi_targets[692] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.half_adder_2.y;
alias fi_targets[693] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.c0;
alias fi_targets[694] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.c1;
alias fi_targets[695] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.ci;
alias fi_targets[696] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.cout;
alias fi_targets[697] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.s;
alias fi_targets[698] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.s0;
alias fi_targets[699] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.x;
alias fi_targets[700] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[17].first_stage.y;
alias fi_targets[701] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.half_adder_1.cout;
alias fi_targets[702] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.half_adder_1.s;
alias fi_targets[703] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.half_adder_1.x;
alias fi_targets[704] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.half_adder_1.y;
alias fi_targets[705] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.half_adder_2.cout;
alias fi_targets[706] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.half_adder_2.s;
alias fi_targets[707] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.half_adder_2.x;
alias fi_targets[708] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.half_adder_2.y;
alias fi_targets[709] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.c0;
alias fi_targets[710] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.c1;
alias fi_targets[711] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.ci;
alias fi_targets[712] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.cout;
alias fi_targets[713] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.s;
alias fi_targets[714] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.s0;
alias fi_targets[715] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.x;
alias fi_targets[716] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[18].first_stage.y;
alias fi_targets[717] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.half_adder_1.cout;
alias fi_targets[718] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.half_adder_1.s;
alias fi_targets[719] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.half_adder_1.x;
alias fi_targets[720] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.half_adder_1.y;
alias fi_targets[721] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.half_adder_2.cout;
alias fi_targets[722] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.half_adder_2.s;
alias fi_targets[723] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.half_adder_2.x;
alias fi_targets[724] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.half_adder_2.y;
alias fi_targets[725] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.c0;
alias fi_targets[726] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.c1;
alias fi_targets[727] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.ci;
alias fi_targets[728] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.cout;
alias fi_targets[729] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.s;
alias fi_targets[730] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.s0;
alias fi_targets[731] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.x;
alias fi_targets[732] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[19].first_stage.y;
alias fi_targets[733] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.half_adder_1.cout;
alias fi_targets[734] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.half_adder_1.s;
alias fi_targets[735] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.half_adder_1.x;
alias fi_targets[736] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.half_adder_1.y;
alias fi_targets[737] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.half_adder_2.cout;
alias fi_targets[738] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.half_adder_2.s;
alias fi_targets[739] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.half_adder_2.x;
alias fi_targets[740] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.half_adder_2.y;
alias fi_targets[741] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.c0;
alias fi_targets[742] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.c1;
alias fi_targets[743] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.ci;
alias fi_targets[744] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.cout;
alias fi_targets[745] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.s;
alias fi_targets[746] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.s0;
alias fi_targets[747] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.x;
alias fi_targets[748] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[1].first_stage.y;
alias fi_targets[749] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.half_adder_1.cout;
alias fi_targets[750] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.half_adder_1.s;
alias fi_targets[751] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.half_adder_1.x;
alias fi_targets[752] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.half_adder_1.y;
alias fi_targets[753] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.half_adder_2.cout;
alias fi_targets[754] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.half_adder_2.s;
alias fi_targets[755] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.half_adder_2.x;
alias fi_targets[756] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.half_adder_2.y;
alias fi_targets[757] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.c0;
alias fi_targets[758] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.c1;
alias fi_targets[759] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.ci;
alias fi_targets[760] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.cout;
alias fi_targets[761] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.s;
alias fi_targets[762] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.s0;
alias fi_targets[763] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.x;
alias fi_targets[764] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[20].first_stage.y;
alias fi_targets[765] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.half_adder_1.cout;
alias fi_targets[766] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.half_adder_1.s;
alias fi_targets[767] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.half_adder_1.x;
alias fi_targets[768] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.half_adder_1.y;
alias fi_targets[769] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.half_adder_2.cout;
alias fi_targets[770] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.half_adder_2.s;
alias fi_targets[771] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.half_adder_2.x;
alias fi_targets[772] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.half_adder_2.y;
alias fi_targets[773] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.c0;
alias fi_targets[774] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.c1;
alias fi_targets[775] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.ci;
alias fi_targets[776] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.cout;
alias fi_targets[777] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.s;
alias fi_targets[778] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.s0;
alias fi_targets[779] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.x;
alias fi_targets[780] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[21].first_stage.y;
alias fi_targets[781] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.half_adder_1.cout;
alias fi_targets[782] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.half_adder_1.s;
alias fi_targets[783] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.half_adder_1.x;
alias fi_targets[784] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.half_adder_1.y;
alias fi_targets[785] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.half_adder_2.cout;
alias fi_targets[786] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.half_adder_2.s;
alias fi_targets[787] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.half_adder_2.x;
alias fi_targets[788] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.half_adder_2.y;
alias fi_targets[789] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.c0;
alias fi_targets[790] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.c1;
alias fi_targets[791] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.ci;
alias fi_targets[792] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.cout;
alias fi_targets[793] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.s;
alias fi_targets[794] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.s0;
alias fi_targets[795] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.x;
alias fi_targets[796] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[22].first_stage.y;
alias fi_targets[797] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.half_adder_1.cout;
alias fi_targets[798] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.half_adder_1.s;
alias fi_targets[799] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.half_adder_1.x;
alias fi_targets[800] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.half_adder_1.y;
alias fi_targets[801] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.half_adder_2.cout;
alias fi_targets[802] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.half_adder_2.s;
alias fi_targets[803] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.half_adder_2.x;
alias fi_targets[804] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.half_adder_2.y;
alias fi_targets[805] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.c0;
alias fi_targets[806] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.c1;
alias fi_targets[807] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.ci;
alias fi_targets[808] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.cout;
alias fi_targets[809] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.s;
alias fi_targets[810] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.s0;
alias fi_targets[811] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.x;
alias fi_targets[812] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[23].first_stage.y;
alias fi_targets[813] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.half_adder_1.cout;
alias fi_targets[814] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.half_adder_1.s;
alias fi_targets[815] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.half_adder_1.x;
alias fi_targets[816] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.half_adder_1.y;
alias fi_targets[817] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.half_adder_2.cout;
alias fi_targets[818] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.half_adder_2.s;
alias fi_targets[819] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.half_adder_2.x;
alias fi_targets[820] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.half_adder_2.y;
alias fi_targets[821] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.c0;
alias fi_targets[822] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.c1;
alias fi_targets[823] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.ci;
alias fi_targets[824] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.cout;
alias fi_targets[825] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.s;
alias fi_targets[826] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.s0;
alias fi_targets[827] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.x;
alias fi_targets[828] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[24].first_stage.y;
alias fi_targets[829] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.half_adder_1.cout;
alias fi_targets[830] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.half_adder_1.s;
alias fi_targets[831] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.half_adder_1.x;
alias fi_targets[832] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.half_adder_1.y;
alias fi_targets[833] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.half_adder_2.cout;
alias fi_targets[834] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.half_adder_2.s;
alias fi_targets[835] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.half_adder_2.x;
alias fi_targets[836] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.half_adder_2.y;
alias fi_targets[837] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.c0;
alias fi_targets[838] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.c1;
alias fi_targets[839] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.ci;
alias fi_targets[840] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.cout;
alias fi_targets[841] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.s;
alias fi_targets[842] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.s0;
alias fi_targets[843] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.x;
alias fi_targets[844] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[25].first_stage.y;
alias fi_targets[845] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.half_adder_1.cout;
alias fi_targets[846] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.half_adder_1.s;
alias fi_targets[847] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.half_adder_1.x;
alias fi_targets[848] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.half_adder_1.y;
alias fi_targets[849] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.half_adder_2.cout;
alias fi_targets[850] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.half_adder_2.s;
alias fi_targets[851] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.half_adder_2.x;
alias fi_targets[852] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.half_adder_2.y;
alias fi_targets[853] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.c0;
alias fi_targets[854] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.c1;
alias fi_targets[855] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.ci;
alias fi_targets[856] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.cout;
alias fi_targets[857] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.s;
alias fi_targets[858] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.s0;
alias fi_targets[859] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.x;
alias fi_targets[860] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[26].first_stage.y;
alias fi_targets[861] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.half_adder_1.cout;
alias fi_targets[862] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.half_adder_1.s;
alias fi_targets[863] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.half_adder_1.x;
alias fi_targets[864] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.half_adder_1.y;
alias fi_targets[865] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.half_adder_2.cout;
alias fi_targets[866] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.half_adder_2.s;
alias fi_targets[867] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.half_adder_2.x;
alias fi_targets[868] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.half_adder_2.y;
alias fi_targets[869] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.c0;
alias fi_targets[870] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.c1;
alias fi_targets[871] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.ci;
alias fi_targets[872] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.cout;
alias fi_targets[873] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.s;
alias fi_targets[874] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.s0;
alias fi_targets[875] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.x;
alias fi_targets[876] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[27].first_stage.y;
alias fi_targets[877] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.half_adder_1.cout;
alias fi_targets[878] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.half_adder_1.s;
alias fi_targets[879] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.half_adder_1.x;
alias fi_targets[880] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.half_adder_1.y;
alias fi_targets[881] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.half_adder_2.cout;
alias fi_targets[882] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.half_adder_2.s;
alias fi_targets[883] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.half_adder_2.x;
alias fi_targets[884] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.half_adder_2.y;
alias fi_targets[885] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.c0;
alias fi_targets[886] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.c1;
alias fi_targets[887] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.ci;
alias fi_targets[888] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.cout;
alias fi_targets[889] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.s;
alias fi_targets[890] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.s0;
alias fi_targets[891] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.x;
alias fi_targets[892] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[28].first_stage.y;
alias fi_targets[893] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.half_adder_1.cout;
alias fi_targets[894] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.half_adder_1.s;
alias fi_targets[895] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.half_adder_1.x;
alias fi_targets[896] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.half_adder_1.y;
alias fi_targets[897] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.half_adder_2.cout;
alias fi_targets[898] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.half_adder_2.s;
alias fi_targets[899] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.half_adder_2.x;
alias fi_targets[900] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.half_adder_2.y;
alias fi_targets[901] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.c0;
alias fi_targets[902] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.c1;
alias fi_targets[903] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.ci;
alias fi_targets[904] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.cout;
alias fi_targets[905] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.s;
alias fi_targets[906] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.s0;
alias fi_targets[907] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.x;
alias fi_targets[908] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[29].first_stage.y;
alias fi_targets[909] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.half_adder_1.cout;
alias fi_targets[910] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.half_adder_1.s;
alias fi_targets[911] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.half_adder_1.x;
alias fi_targets[912] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.half_adder_1.y;
alias fi_targets[913] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.half_adder_2.cout;
alias fi_targets[914] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.half_adder_2.s;
alias fi_targets[915] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.half_adder_2.x;
alias fi_targets[916] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.half_adder_2.y;
alias fi_targets[917] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.c0;
alias fi_targets[918] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.c1;
alias fi_targets[919] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.ci;
alias fi_targets[920] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.cout;
alias fi_targets[921] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.s;
alias fi_targets[922] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.s0;
alias fi_targets[923] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.x;
alias fi_targets[924] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[2].first_stage.y;
alias fi_targets[925] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.half_adder_1.cout;
alias fi_targets[926] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.half_adder_1.s;
alias fi_targets[927] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.half_adder_1.x;
alias fi_targets[928] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.half_adder_1.y;
alias fi_targets[929] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.half_adder_2.cout;
alias fi_targets[930] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.half_adder_2.s;
alias fi_targets[931] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.half_adder_2.x;
alias fi_targets[932] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.half_adder_2.y;
alias fi_targets[933] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.c0;
alias fi_targets[934] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.c1;
alias fi_targets[935] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.ci;
alias fi_targets[936] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.cout;
alias fi_targets[937] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.s;
alias fi_targets[938] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.s0;
alias fi_targets[939] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.x;
alias fi_targets[940] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[30].first_stage.y;
alias fi_targets[941] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.half_adder_1.cout;
alias fi_targets[942] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.half_adder_1.s;
alias fi_targets[943] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.half_adder_1.x;
alias fi_targets[944] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.half_adder_1.y;
alias fi_targets[945] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.half_adder_2.cout;
alias fi_targets[946] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.half_adder_2.s;
alias fi_targets[947] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.half_adder_2.x;
alias fi_targets[948] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.half_adder_2.y;
alias fi_targets[949] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.c0;
alias fi_targets[950] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.c1;
alias fi_targets[951] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.ci;
alias fi_targets[952] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.cout;
alias fi_targets[953] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.s;
alias fi_targets[954] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.s0;
alias fi_targets[955] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.x;
alias fi_targets[956] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[31].first_stage.y;
alias fi_targets[957] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.half_adder_1.cout;
alias fi_targets[958] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.half_adder_1.s;
alias fi_targets[959] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.half_adder_1.x;
alias fi_targets[960] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.half_adder_1.y;
alias fi_targets[961] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.half_adder_2.cout;
alias fi_targets[962] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.half_adder_2.s;
alias fi_targets[963] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.half_adder_2.x;
alias fi_targets[964] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.half_adder_2.y;
alias fi_targets[965] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.c0;
alias fi_targets[966] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.c1;
alias fi_targets[967] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.ci;
alias fi_targets[968] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.cout;
alias fi_targets[969] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.s;
alias fi_targets[970] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.s0;
alias fi_targets[971] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.x;
alias fi_targets[972] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[3].first_stage.y;
alias fi_targets[973] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.half_adder_1.cout;
alias fi_targets[974] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.half_adder_1.s;
alias fi_targets[975] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.half_adder_1.x;
alias fi_targets[976] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.half_adder_1.y;
alias fi_targets[977] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.half_adder_2.cout;
alias fi_targets[978] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.half_adder_2.s;
alias fi_targets[979] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.half_adder_2.x;
alias fi_targets[980] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.half_adder_2.y;
alias fi_targets[981] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.c0;
alias fi_targets[982] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.c1;
alias fi_targets[983] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.ci;
alias fi_targets[984] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.cout;
alias fi_targets[985] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.s;
alias fi_targets[986] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.s0;
alias fi_targets[987] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.x;
alias fi_targets[988] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[4].first_stage.y;
alias fi_targets[989] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.half_adder_1.cout;
alias fi_targets[990] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.half_adder_1.s;
alias fi_targets[991] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.half_adder_1.x;
alias fi_targets[992] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.half_adder_1.y;
alias fi_targets[993] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.half_adder_2.cout;
alias fi_targets[994] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.half_adder_2.s;
alias fi_targets[995] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.half_adder_2.x;
alias fi_targets[996] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.half_adder_2.y;
alias fi_targets[997] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.c0;
alias fi_targets[998] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.c1;
alias fi_targets[999] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.ci;
alias fi_targets[1000] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.cout;
alias fi_targets[1001] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.s;
alias fi_targets[1002] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.s0;
alias fi_targets[1003] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.x;
alias fi_targets[1004] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[5].first_stage.y;
alias fi_targets[1005] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.half_adder_1.cout;
alias fi_targets[1006] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.half_adder_1.s;
alias fi_targets[1007] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.half_adder_1.x;
alias fi_targets[1008] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.half_adder_1.y;
alias fi_targets[1009] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.half_adder_2.cout;
alias fi_targets[1010] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.half_adder_2.s;
alias fi_targets[1011] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.half_adder_2.x;
alias fi_targets[1012] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.half_adder_2.y;
alias fi_targets[1013] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.c0;
alias fi_targets[1014] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.c1;
alias fi_targets[1015] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.ci;
alias fi_targets[1016] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.cout;
alias fi_targets[1017] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.s;
alias fi_targets[1018] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.s0;
alias fi_targets[1019] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.x;
alias fi_targets[1020] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[6].first_stage.y;
alias fi_targets[1021] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.half_adder_1.cout;
alias fi_targets[1022] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.half_adder_1.s;
alias fi_targets[1023] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.half_adder_1.x;
alias fi_targets[1024] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.half_adder_1.y;
alias fi_targets[1025] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.half_adder_2.cout;
alias fi_targets[1026] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.half_adder_2.s;
alias fi_targets[1027] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.half_adder_2.x;
alias fi_targets[1028] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.half_adder_2.y;
alias fi_targets[1029] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.c0;
alias fi_targets[1030] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.c1;
alias fi_targets[1031] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.ci;
alias fi_targets[1032] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.cout;
alias fi_targets[1033] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.s;
alias fi_targets[1034] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.s0;
alias fi_targets[1035] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.x;
alias fi_targets[1036] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[7].first_stage.y;
alias fi_targets[1037] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.half_adder_1.cout;
alias fi_targets[1038] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.half_adder_1.s;
alias fi_targets[1039] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.half_adder_1.x;
alias fi_targets[1040] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.half_adder_1.y;
alias fi_targets[1041] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.half_adder_2.cout;
alias fi_targets[1042] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.half_adder_2.s;
alias fi_targets[1043] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.half_adder_2.x;
alias fi_targets[1044] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.half_adder_2.y;
alias fi_targets[1045] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.c0;
alias fi_targets[1046] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.c1;
alias fi_targets[1047] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.ci;
alias fi_targets[1048] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.cout;
alias fi_targets[1049] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.s;
alias fi_targets[1050] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.s0;
alias fi_targets[1051] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.x;
alias fi_targets[1052] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[8].first_stage.y;
alias fi_targets[1053] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.half_adder_1.cout;
alias fi_targets[1054] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.half_adder_1.s;
alias fi_targets[1055] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.half_adder_1.x;
alias fi_targets[1056] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.half_adder_1.y;
alias fi_targets[1057] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.half_adder_2.cout;
alias fi_targets[1058] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.half_adder_2.s;
alias fi_targets[1059] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.half_adder_2.x;
alias fi_targets[1060] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.half_adder_2.y;
alias fi_targets[1061] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.c0;
alias fi_targets[1062] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.c1;
alias fi_targets[1063] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.ci;
alias fi_targets[1064] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.cout;
alias fi_targets[1065] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.s;
alias fi_targets[1066] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.s0;
alias fi_targets[1067] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.x;
alias fi_targets[1068] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.genblk1[9].first_stage.y;
alias fi_targets[1069] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.A;
alias fi_targets[1070] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.B;
alias fi_targets[1071] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.C;
alias fi_targets[1072] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.C1;
alias fi_targets[1073] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.RCA_out;
alias fi_targets[1074] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.S;
alias fi_targets[1075] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.S1;
alias fi_targets[1076] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.cout;
alias fi_targets[1077] = dv_top.dut.EX.func_unit.alu.arithmetic.ADD_SUB.v;
alias fi_targets[1078] = dv_top.dut.EX.func_unit.alu.arithmetic.n_mux.addr;
alias fi_targets[1079] = dv_top.dut.EX.func_unit.alu.arithmetic.n_mux.data_in;
alias fi_targets[1080] = dv_top.dut.EX.func_unit.alu.arithmetic.n_mux.data_out;
alias fi_targets[1081] = dv_top.dut.EX.func_unit.alu.arithmetic.n_mux.inner_data;
alias fi_targets[1082] = dv_top.dut.EX.func_unit.alu.arithmetic.out_mux.addr;
alias fi_targets[1083] = dv_top.dut.EX.func_unit.alu.arithmetic.out_mux.data_in;
alias fi_targets[1084] = dv_top.dut.EX.func_unit.alu.arithmetic.out_mux.data_out;
alias fi_targets[1085] = dv_top.dut.EX.func_unit.alu.arithmetic.out_mux.inner_data;
alias fi_targets[1086] = dv_top.dut.EX.func_unit.alu.arithmetic.add_sub_out;
alias fi_targets[1087] = dv_top.dut.EX.func_unit.alu.arithmetic.carry_out;
alias fi_targets[1088] = dv_top.dut.EX.func_unit.alu.arithmetic.data_a;
alias fi_targets[1089] = dv_top.dut.EX.func_unit.alu.arithmetic.data_b;
alias fi_targets[1090] = dv_top.dut.EX.func_unit.alu.arithmetic.data_b_prep;
alias fi_targets[1091] = dv_top.dut.EX.func_unit.alu.arithmetic.data_result;
alias fi_targets[1092] = dv_top.dut.EX.func_unit.alu.arithmetic.func_sel;
alias fi_targets[1093] = dv_top.dut.EX.func_unit.alu.arithmetic.negative;
alias fi_targets[1094] = dv_top.dut.EX.func_unit.alu.arithmetic.out_select;
alias fi_targets[1095] = dv_top.dut.EX.func_unit.alu.arithmetic.overflow;
alias fi_targets[1096] = dv_top.dut.EX.func_unit.alu.arithmetic.sub;
alias fi_targets[1097] = dv_top.dut.EX.func_unit.alu.arithmetic.usign;
alias fi_targets[1098] = dv_top.dut.EX.func_unit.alu.arithmetic.zero;
alias fi_targets[1099] = dv_top.dut.EX.func_unit.alu.logical.out_mux.addr;
alias fi_targets[1100] = dv_top.dut.EX.func_unit.alu.logical.out_mux.data_in;
alias fi_targets[1101] = dv_top.dut.EX.func_unit.alu.logical.out_mux.data_out;
alias fi_targets[1102] = dv_top.dut.EX.func_unit.alu.logical.out_mux.inner_data;
alias fi_targets[1103] = dv_top.dut.EX.func_unit.alu.logical.and_result;
alias fi_targets[1104] = dv_top.dut.EX.func_unit.alu.logical.data_a;
alias fi_targets[1105] = dv_top.dut.EX.func_unit.alu.logical.data_b;
alias fi_targets[1106] = dv_top.dut.EX.func_unit.alu.logical.data_result;
alias fi_targets[1107] = dv_top.dut.EX.func_unit.alu.logical.func_sel;
alias fi_targets[1108] = dv_top.dut.EX.func_unit.alu.logical.or_result;
alias fi_targets[1109] = dv_top.dut.EX.func_unit.alu.logical.xor_result;
alias fi_targets[1110] = dv_top.dut.EX.func_unit.alu.out_mux.addr;
alias fi_targets[1111] = dv_top.dut.EX.func_unit.alu.out_mux.data_in;
alias fi_targets[1112] = dv_top.dut.EX.func_unit.alu.out_mux.data_out;
alias fi_targets[1113] = dv_top.dut.EX.func_unit.alu.out_mux.inner_data;
alias fi_targets[1114] = dv_top.dut.EX.func_unit.alu.arithmetic_out;
alias fi_targets[1115] = dv_top.dut.EX.func_unit.alu.carry_out;
alias fi_targets[1116] = dv_top.dut.EX.func_unit.alu.data_a;
alias fi_targets[1117] = dv_top.dut.EX.func_unit.alu.data_b;
alias fi_targets[1118] = dv_top.dut.EX.func_unit.alu.data_result;
alias fi_targets[1119] = dv_top.dut.EX.func_unit.alu.func_sel;
alias fi_targets[1120] = dv_top.dut.EX.func_unit.alu.logical_out;
alias fi_targets[1121] = dv_top.dut.EX.func_unit.alu.negative;
alias fi_targets[1122] = dv_top.dut.EX.func_unit.alu.overflow;
alias fi_targets[1123] = dv_top.dut.EX.func_unit.alu.zero;
alias fi_targets[1124] = dv_top.dut.EX.func_unit.out_mux.addr;
alias fi_targets[1125] = dv_top.dut.EX.func_unit.out_mux.data_in;
alias fi_targets[1126] = dv_top.dut.EX.func_unit.out_mux.data_out;
alias fi_targets[1127] = dv_top.dut.EX.func_unit.out_mux.inner_data;
alias fi_targets[1128] = dv_top.dut.EX.func_unit.shifter.genblk2[0].mux.addr;
alias fi_targets[1129] = dv_top.dut.EX.func_unit.shifter.genblk2[0].mux.data_in;
alias fi_targets[1130] = dv_top.dut.EX.func_unit.shifter.genblk2[0].mux.data_out;
alias fi_targets[1131] = dv_top.dut.EX.func_unit.shifter.genblk2[0].mux.inner_data;
alias fi_targets[1132] = dv_top.dut.EX.func_unit.shifter.genblk2[10].mux.addr;
alias fi_targets[1133] = dv_top.dut.EX.func_unit.shifter.genblk2[10].mux.data_in;
alias fi_targets[1134] = dv_top.dut.EX.func_unit.shifter.genblk2[10].mux.data_out;
alias fi_targets[1135] = dv_top.dut.EX.func_unit.shifter.genblk2[10].mux.inner_data;
alias fi_targets[1136] = dv_top.dut.EX.func_unit.shifter.genblk2[11].mux.addr;
alias fi_targets[1137] = dv_top.dut.EX.func_unit.shifter.genblk2[11].mux.data_in;
alias fi_targets[1138] = dv_top.dut.EX.func_unit.shifter.genblk2[11].mux.data_out;
alias fi_targets[1139] = dv_top.dut.EX.func_unit.shifter.genblk2[11].mux.inner_data;
alias fi_targets[1140] = dv_top.dut.EX.func_unit.shifter.genblk2[12].mux.addr;
alias fi_targets[1141] = dv_top.dut.EX.func_unit.shifter.genblk2[12].mux.data_in;
alias fi_targets[1142] = dv_top.dut.EX.func_unit.shifter.genblk2[12].mux.data_out;
alias fi_targets[1143] = dv_top.dut.EX.func_unit.shifter.genblk2[12].mux.inner_data;
alias fi_targets[1144] = dv_top.dut.EX.func_unit.shifter.genblk2[13].mux.addr;
alias fi_targets[1145] = dv_top.dut.EX.func_unit.shifter.genblk2[13].mux.data_in;
alias fi_targets[1146] = dv_top.dut.EX.func_unit.shifter.genblk2[13].mux.data_out;
alias fi_targets[1147] = dv_top.dut.EX.func_unit.shifter.genblk2[13].mux.inner_data;
alias fi_targets[1148] = dv_top.dut.EX.func_unit.shifter.genblk2[14].mux.addr;
alias fi_targets[1149] = dv_top.dut.EX.func_unit.shifter.genblk2[14].mux.data_in;
alias fi_targets[1150] = dv_top.dut.EX.func_unit.shifter.genblk2[14].mux.data_out;
alias fi_targets[1151] = dv_top.dut.EX.func_unit.shifter.genblk2[14].mux.inner_data;
alias fi_targets[1152] = dv_top.dut.EX.func_unit.shifter.genblk2[15].mux.addr;
alias fi_targets[1153] = dv_top.dut.EX.func_unit.shifter.genblk2[15].mux.data_in;
alias fi_targets[1154] = dv_top.dut.EX.func_unit.shifter.genblk2[15].mux.data_out;
alias fi_targets[1155] = dv_top.dut.EX.func_unit.shifter.genblk2[15].mux.inner_data;
alias fi_targets[1156] = dv_top.dut.EX.func_unit.shifter.genblk2[16].mux.addr;
alias fi_targets[1157] = dv_top.dut.EX.func_unit.shifter.genblk2[16].mux.data_in;
alias fi_targets[1158] = dv_top.dut.EX.func_unit.shifter.genblk2[16].mux.data_out;
alias fi_targets[1159] = dv_top.dut.EX.func_unit.shifter.genblk2[16].mux.inner_data;
alias fi_targets[1160] = dv_top.dut.EX.func_unit.shifter.genblk2[17].mux.addr;
alias fi_targets[1161] = dv_top.dut.EX.func_unit.shifter.genblk2[17].mux.data_in;
alias fi_targets[1162] = dv_top.dut.EX.func_unit.shifter.genblk2[17].mux.data_out;
alias fi_targets[1163] = dv_top.dut.EX.func_unit.shifter.genblk2[17].mux.inner_data;
alias fi_targets[1164] = dv_top.dut.EX.func_unit.shifter.genblk2[18].mux.addr;
alias fi_targets[1165] = dv_top.dut.EX.func_unit.shifter.genblk2[18].mux.data_in;
alias fi_targets[1166] = dv_top.dut.EX.func_unit.shifter.genblk2[18].mux.data_out;
alias fi_targets[1167] = dv_top.dut.EX.func_unit.shifter.genblk2[18].mux.inner_data;
alias fi_targets[1168] = dv_top.dut.EX.func_unit.shifter.genblk2[19].mux.addr;
alias fi_targets[1169] = dv_top.dut.EX.func_unit.shifter.genblk2[19].mux.data_in;
alias fi_targets[1170] = dv_top.dut.EX.func_unit.shifter.genblk2[19].mux.data_out;
alias fi_targets[1171] = dv_top.dut.EX.func_unit.shifter.genblk2[19].mux.inner_data;
alias fi_targets[1172] = dv_top.dut.EX.func_unit.shifter.genblk2[1].mux.addr;
alias fi_targets[1173] = dv_top.dut.EX.func_unit.shifter.genblk2[1].mux.data_in;
alias fi_targets[1174] = dv_top.dut.EX.func_unit.shifter.genblk2[1].mux.data_out;
alias fi_targets[1175] = dv_top.dut.EX.func_unit.shifter.genblk2[1].mux.inner_data;
alias fi_targets[1176] = dv_top.dut.EX.func_unit.shifter.genblk2[20].mux.addr;
alias fi_targets[1177] = dv_top.dut.EX.func_unit.shifter.genblk2[20].mux.data_in;
alias fi_targets[1178] = dv_top.dut.EX.func_unit.shifter.genblk2[20].mux.data_out;
alias fi_targets[1179] = dv_top.dut.EX.func_unit.shifter.genblk2[20].mux.inner_data;
alias fi_targets[1180] = dv_top.dut.EX.func_unit.shifter.genblk2[21].mux.addr;
alias fi_targets[1181] = dv_top.dut.EX.func_unit.shifter.genblk2[21].mux.data_in;
alias fi_targets[1182] = dv_top.dut.EX.func_unit.shifter.genblk2[21].mux.data_out;
alias fi_targets[1183] = dv_top.dut.EX.func_unit.shifter.genblk2[21].mux.inner_data;
alias fi_targets[1184] = dv_top.dut.EX.func_unit.shifter.genblk2[22].mux.addr;
alias fi_targets[1185] = dv_top.dut.EX.func_unit.shifter.genblk2[22].mux.data_in;
alias fi_targets[1186] = dv_top.dut.EX.func_unit.shifter.genblk2[22].mux.data_out;
alias fi_targets[1187] = dv_top.dut.EX.func_unit.shifter.genblk2[22].mux.inner_data;
alias fi_targets[1188] = dv_top.dut.EX.func_unit.shifter.genblk2[23].mux.addr;
alias fi_targets[1189] = dv_top.dut.EX.func_unit.shifter.genblk2[23].mux.data_in;
alias fi_targets[1190] = dv_top.dut.EX.func_unit.shifter.genblk2[23].mux.data_out;
alias fi_targets[1191] = dv_top.dut.EX.func_unit.shifter.genblk2[23].mux.inner_data;
alias fi_targets[1192] = dv_top.dut.EX.func_unit.shifter.genblk2[24].mux.addr;
alias fi_targets[1193] = dv_top.dut.EX.func_unit.shifter.genblk2[24].mux.data_in;
alias fi_targets[1194] = dv_top.dut.EX.func_unit.shifter.genblk2[24].mux.data_out;
alias fi_targets[1195] = dv_top.dut.EX.func_unit.shifter.genblk2[24].mux.inner_data;
alias fi_targets[1196] = dv_top.dut.EX.func_unit.shifter.genblk2[25].mux.addr;
alias fi_targets[1197] = dv_top.dut.EX.func_unit.shifter.genblk2[25].mux.data_in;
alias fi_targets[1198] = dv_top.dut.EX.func_unit.shifter.genblk2[25].mux.data_out;
alias fi_targets[1199] = dv_top.dut.EX.func_unit.shifter.genblk2[25].mux.inner_data;
alias fi_targets[1200] = dv_top.dut.EX.func_unit.shifter.genblk2[26].mux.addr;
alias fi_targets[1201] = dv_top.dut.EX.func_unit.shifter.genblk2[26].mux.data_in;
alias fi_targets[1202] = dv_top.dut.EX.func_unit.shifter.genblk2[26].mux.data_out;
alias fi_targets[1203] = dv_top.dut.EX.func_unit.shifter.genblk2[26].mux.inner_data;
alias fi_targets[1204] = dv_top.dut.EX.func_unit.shifter.genblk2[27].mux.addr;
alias fi_targets[1205] = dv_top.dut.EX.func_unit.shifter.genblk2[27].mux.data_in;
alias fi_targets[1206] = dv_top.dut.EX.func_unit.shifter.genblk2[27].mux.data_out;
alias fi_targets[1207] = dv_top.dut.EX.func_unit.shifter.genblk2[27].mux.inner_data;
alias fi_targets[1208] = dv_top.dut.EX.func_unit.shifter.genblk2[28].mux.addr;
alias fi_targets[1209] = dv_top.dut.EX.func_unit.shifter.genblk2[28].mux.data_in;
alias fi_targets[1210] = dv_top.dut.EX.func_unit.shifter.genblk2[28].mux.data_out;
alias fi_targets[1211] = dv_top.dut.EX.func_unit.shifter.genblk2[28].mux.inner_data;
alias fi_targets[1212] = dv_top.dut.EX.func_unit.shifter.genblk2[29].mux.addr;
alias fi_targets[1213] = dv_top.dut.EX.func_unit.shifter.genblk2[29].mux.data_in;
alias fi_targets[1214] = dv_top.dut.EX.func_unit.shifter.genblk2[29].mux.data_out;
alias fi_targets[1215] = dv_top.dut.EX.func_unit.shifter.genblk2[29].mux.inner_data;
alias fi_targets[1216] = dv_top.dut.EX.func_unit.shifter.genblk2[2].mux.addr;
alias fi_targets[1217] = dv_top.dut.EX.func_unit.shifter.genblk2[2].mux.data_in;
alias fi_targets[1218] = dv_top.dut.EX.func_unit.shifter.genblk2[2].mux.data_out;
alias fi_targets[1219] = dv_top.dut.EX.func_unit.shifter.genblk2[2].mux.inner_data;
alias fi_targets[1220] = dv_top.dut.EX.func_unit.shifter.genblk2[30].mux.addr;
alias fi_targets[1221] = dv_top.dut.EX.func_unit.shifter.genblk2[30].mux.data_in;
alias fi_targets[1222] = dv_top.dut.EX.func_unit.shifter.genblk2[30].mux.data_out;
alias fi_targets[1223] = dv_top.dut.EX.func_unit.shifter.genblk2[30].mux.inner_data;
alias fi_targets[1224] = dv_top.dut.EX.func_unit.shifter.genblk2[31].mux.addr;
alias fi_targets[1225] = dv_top.dut.EX.func_unit.shifter.genblk2[31].mux.data_in;
alias fi_targets[1226] = dv_top.dut.EX.func_unit.shifter.genblk2[31].mux.data_out;
alias fi_targets[1227] = dv_top.dut.EX.func_unit.shifter.genblk2[31].mux.inner_data;
alias fi_targets[1228] = dv_top.dut.EX.func_unit.shifter.genblk2[3].mux.addr;
alias fi_targets[1229] = dv_top.dut.EX.func_unit.shifter.genblk2[3].mux.data_in;
alias fi_targets[1230] = dv_top.dut.EX.func_unit.shifter.genblk2[3].mux.data_out;
alias fi_targets[1231] = dv_top.dut.EX.func_unit.shifter.genblk2[3].mux.inner_data;
alias fi_targets[1232] = dv_top.dut.EX.func_unit.shifter.genblk2[4].mux.addr;
alias fi_targets[1233] = dv_top.dut.EX.func_unit.shifter.genblk2[4].mux.data_in;
alias fi_targets[1234] = dv_top.dut.EX.func_unit.shifter.genblk2[4].mux.data_out;
alias fi_targets[1235] = dv_top.dut.EX.func_unit.shifter.genblk2[4].mux.inner_data;
alias fi_targets[1236] = dv_top.dut.EX.func_unit.shifter.genblk2[5].mux.addr;
alias fi_targets[1237] = dv_top.dut.EX.func_unit.shifter.genblk2[5].mux.data_in;
alias fi_targets[1238] = dv_top.dut.EX.func_unit.shifter.genblk2[5].mux.data_out;
alias fi_targets[1239] = dv_top.dut.EX.func_unit.shifter.genblk2[5].mux.inner_data;
alias fi_targets[1240] = dv_top.dut.EX.func_unit.shifter.genblk2[6].mux.addr;
alias fi_targets[1241] = dv_top.dut.EX.func_unit.shifter.genblk2[6].mux.data_in;
alias fi_targets[1242] = dv_top.dut.EX.func_unit.shifter.genblk2[6].mux.data_out;
alias fi_targets[1243] = dv_top.dut.EX.func_unit.shifter.genblk2[6].mux.inner_data;
alias fi_targets[1244] = dv_top.dut.EX.func_unit.shifter.genblk2[7].mux.addr;
alias fi_targets[1245] = dv_top.dut.EX.func_unit.shifter.genblk2[7].mux.data_in;
alias fi_targets[1246] = dv_top.dut.EX.func_unit.shifter.genblk2[7].mux.data_out;
alias fi_targets[1247] = dv_top.dut.EX.func_unit.shifter.genblk2[7].mux.inner_data;
alias fi_targets[1248] = dv_top.dut.EX.func_unit.shifter.genblk2[8].mux.addr;
alias fi_targets[1249] = dv_top.dut.EX.func_unit.shifter.genblk2[8].mux.data_in;
alias fi_targets[1250] = dv_top.dut.EX.func_unit.shifter.genblk2[8].mux.data_out;
alias fi_targets[1251] = dv_top.dut.EX.func_unit.shifter.genblk2[8].mux.inner_data;
alias fi_targets[1252] = dv_top.dut.EX.func_unit.shifter.genblk2[9].mux.addr;
alias fi_targets[1253] = dv_top.dut.EX.func_unit.shifter.genblk2[9].mux.data_in;
alias fi_targets[1254] = dv_top.dut.EX.func_unit.shifter.genblk2[9].mux.data_out;
alias fi_targets[1255] = dv_top.dut.EX.func_unit.shifter.genblk2[9].mux.inner_data;
alias fi_targets[1256] = dv_top.dut.EX.func_unit.shifter.Data_in;
alias fi_targets[1257] = dv_top.dut.EX.func_unit.shifter.Data_out;
alias fi_targets[1258] = dv_top.dut.EX.func_unit.shifter.Sel;
alias fi_targets[1259] = dv_top.dut.EX.func_unit.shifter.arithmetic_shifter_in;
alias fi_targets[1260] = dv_top.dut.EX.func_unit.shifter.left;
alias fi_targets[1261] = dv_top.dut.EX.func_unit.shifter.shamt;
alias fi_targets[1262] = dv_top.dut.EX.func_unit.shifter.shifter_in;
alias fi_targets[1263] = dv_top.dut.EX.func_unit.shifter.shifter_out;
alias fi_targets[1264] = dv_top.dut.EX.func_unit.alu_c;
alias fi_targets[1265] = dv_top.dut.EX.func_unit.alu_n;
alias fi_targets[1266] = dv_top.dut.EX.func_unit.alu_out;
alias fi_targets[1267] = dv_top.dut.EX.func_unit.alu_v;
alias fi_targets[1268] = dv_top.dut.EX.func_unit.alu_z;
alias fi_targets[1269] = dv_top.dut.EX.func_unit.carry_out;
alias fi_targets[1270] = dv_top.dut.EX.func_unit.data_a;
alias fi_targets[1271] = dv_top.dut.EX.func_unit.data_b;
alias fi_targets[1272] = dv_top.dut.EX.func_unit.data_result;
alias fi_targets[1273] = dv_top.dut.EX.func_unit.func_sel;
alias fi_targets[1274] = dv_top.dut.EX.func_unit.negative;
alias fi_targets[1275] = dv_top.dut.EX.func_unit.overflow;
alias fi_targets[1276] = dv_top.dut.EX.func_unit.shifter_out;
alias fi_targets[1277] = dv_top.dut.EX.func_unit.zero;
alias fi_targets[1278] = dv_top.dut.EX.pc_correction_mux.addr;
alias fi_targets[1279] = dv_top.dut.EX.pc_correction_mux.data_in;
alias fi_targets[1280] = dv_top.dut.EX.pc_correction_mux.data_out;
alias fi_targets[1281] = dv_top.dut.EX.pc_correction_mux.inner_data;
alias fi_targets[1282] = dv_top.dut.EX.pc_mux.addr;
alias fi_targets[1283] = dv_top.dut.EX.pc_mux.data_in;
alias fi_targets[1284] = dv_top.dut.EX.pc_mux.data_out;
alias fi_targets[1285] = dv_top.dut.EX.pc_mux.inner_data;
alias fi_targets[1286] = dv_top.dut.EX.N;
alias fi_targets[1287] = dv_top.dut.EX.Real_MPC;
alias fi_targets[1288] = dv_top.dut.EX.Z;
alias fi_targets[1289] = dv_top.dut.EX.branch_prediction_i;
alias fi_targets[1290] = dv_top.dut.EX.branch_sel;
alias fi_targets[1291] = dv_top.dut.EX.calculated_result_internal;
alias fi_targets[1292] = dv_top.dut.EX.calculated_result_o;
alias fi_targets[1293] = dv_top.dut.EX.control_signal_i;
alias fi_targets[1294] = dv_top.dut.EX.control_signal_internal;
alias fi_targets[1295] = dv_top.dut.EX.control_signal_o;
alias fi_targets[1296] = dv_top.dut.EX.correct_pc;
alias fi_targets[1297] = dv_top.dut.EX.data_a;
alias fi_targets[1298] = dv_top.dut.EX.data_a_forward_sel;
alias fi_targets[1299] = dv_top.dut.EX.data_a_i;
alias fi_targets[1300] = dv_top.dut.EX.data_b;
alias fi_targets[1301] = dv_top.dut.EX.data_b_forward_sel;
alias fi_targets[1302] = dv_top.dut.EX.data_b_i;
alias fi_targets[1303] = dv_top.dut.EX.data_from_mem;
alias fi_targets[1304] = dv_top.dut.EX.data_from_wb;
alias fi_targets[1305] = dv_top.dut.EX.data_store_forward_sel;
alias fi_targets[1306] = dv_top.dut.EX.function_unit_o;
alias fi_targets[1307] = dv_top.dut.EX.isJALR;
alias fi_targets[1308] = dv_top.dut.EX.misprediction_o;
alias fi_targets[1309] = dv_top.dut.EX.pc_plus_i;
alias fi_targets[1310] = dv_top.dut.EX.rs1_addr;
alias fi_targets[1311] = dv_top.dut.EX.rs2_addr;
alias fi_targets[1312] = dv_top.dut.EX.store_data_i;
alias fi_targets[1313] = dv_top.dut.EX.store_data_internal;
alias fi_targets[1314] = dv_top.dut.EX.store_data_o;
alias fi_targets[1315] = dv_top.dut.HD.RA_ID;
alias fi_targets[1316] = dv_top.dut.HD.RB_ID;
alias fi_targets[1317] = dv_top.dut.HD.RD_EX;
alias fi_targets[1318] = dv_top.dut.HD.RD_RA;
alias fi_targets[1319] = dv_top.dut.HD.RD_RB;
alias fi_targets[1320] = dv_top.dut.HD.buble;
alias fi_targets[1321] = dv_top.dut.HD.isLoad_EX;
alias fi_targets[1322] = dv_top.dut.HD.isRA;
alias fi_targets[1323] = dv_top.dut.HD.isRB;
alias fi_targets[1324] = dv_top.dut.ID.Mux_B.addr;
alias fi_targets[1325] = dv_top.dut.ID.Mux_B.data_in;
alias fi_targets[1326] = dv_top.dut.ID.Mux_B.data_out;
alias fi_targets[1327] = dv_top.dut.ID.Mux_B.inner_data;
alias fi_targets[1328] = dv_top.dut.ID.RegFile.a_mux_out.addr;
alias fi_targets[1329] = dv_top.dut.ID.RegFile.a_mux_out.data_in;
alias fi_targets[1330] = dv_top.dut.ID.RegFile.a_mux_out.data_out;
alias fi_targets[1331] = dv_top.dut.ID.RegFile.a_mux_out.inner_data;
alias fi_targets[1332] = dv_top.dut.ID.RegFile.b_mux_out.addr;
alias fi_targets[1333] = dv_top.dut.ID.RegFile.b_mux_out.data_in;
alias fi_targets[1334] = dv_top.dut.ID.RegFile.b_mux_out.data_out;
alias fi_targets[1335] = dv_top.dut.ID.RegFile.b_mux_out.inner_data;
alias fi_targets[1336] = dv_top.dut.ID.RegFile.decoder_in.addr;
alias fi_targets[1337] = dv_top.dut.ID.RegFile.decoder_in.dec_out;
alias fi_targets[1338] = dv_top.dut.ID.RegFile.registers.a0.data_in;
alias fi_targets[1339] = dv_top.dut.ID.RegFile.registers.a0.data_out;
alias fi_targets[1340] = dv_top.dut.ID.RegFile.registers.a0.we;
alias fi_targets[1341] = dv_top.dut.ID.RegFile.registers.a1.data_in;
alias fi_targets[1342] = dv_top.dut.ID.RegFile.registers.a1.data_out;
alias fi_targets[1343] = dv_top.dut.ID.RegFile.registers.a1.we;
alias fi_targets[1344] = dv_top.dut.ID.RegFile.registers.a2.data_in;
alias fi_targets[1345] = dv_top.dut.ID.RegFile.registers.a2.data_out;
alias fi_targets[1346] = dv_top.dut.ID.RegFile.registers.a2.we;
alias fi_targets[1347] = dv_top.dut.ID.RegFile.registers.a3.data_in;
alias fi_targets[1348] = dv_top.dut.ID.RegFile.registers.a3.data_out;
alias fi_targets[1349] = dv_top.dut.ID.RegFile.registers.a3.we;
alias fi_targets[1350] = dv_top.dut.ID.RegFile.registers.a4.data_in;
alias fi_targets[1351] = dv_top.dut.ID.RegFile.registers.a4.data_out;
alias fi_targets[1352] = dv_top.dut.ID.RegFile.registers.a4.we;
alias fi_targets[1353] = dv_top.dut.ID.RegFile.registers.a5.data_in;
alias fi_targets[1354] = dv_top.dut.ID.RegFile.registers.a5.data_out;
alias fi_targets[1355] = dv_top.dut.ID.RegFile.registers.a5.we;
alias fi_targets[1356] = dv_top.dut.ID.RegFile.registers.a6.data_in;
alias fi_targets[1357] = dv_top.dut.ID.RegFile.registers.a6.data_out;
alias fi_targets[1358] = dv_top.dut.ID.RegFile.registers.a6.we;
alias fi_targets[1359] = dv_top.dut.ID.RegFile.registers.a7.data_in;
alias fi_targets[1360] = dv_top.dut.ID.RegFile.registers.a7.data_out;
alias fi_targets[1361] = dv_top.dut.ID.RegFile.registers.a7.we;
alias fi_targets[1362] = dv_top.dut.ID.RegFile.registers.gp.data_in;
alias fi_targets[1363] = dv_top.dut.ID.RegFile.registers.gp.data_out;
alias fi_targets[1364] = dv_top.dut.ID.RegFile.registers.gp.we;
alias fi_targets[1365] = dv_top.dut.ID.RegFile.registers.ra.data_in;
alias fi_targets[1366] = dv_top.dut.ID.RegFile.registers.ra.data_out;
alias fi_targets[1367] = dv_top.dut.ID.RegFile.registers.ra.we;
alias fi_targets[1368] = dv_top.dut.ID.RegFile.registers.s0.data_in;
alias fi_targets[1369] = dv_top.dut.ID.RegFile.registers.s0.data_out;
alias fi_targets[1370] = dv_top.dut.ID.RegFile.registers.s0.we;
alias fi_targets[1371] = dv_top.dut.ID.RegFile.registers.s1.data_in;
alias fi_targets[1372] = dv_top.dut.ID.RegFile.registers.s1.data_out;
alias fi_targets[1373] = dv_top.dut.ID.RegFile.registers.s1.we;
alias fi_targets[1374] = dv_top.dut.ID.RegFile.registers.s10.data_in;
alias fi_targets[1375] = dv_top.dut.ID.RegFile.registers.s10.data_out;
alias fi_targets[1376] = dv_top.dut.ID.RegFile.registers.s10.we;
alias fi_targets[1377] = dv_top.dut.ID.RegFile.registers.s11.data_in;
alias fi_targets[1378] = dv_top.dut.ID.RegFile.registers.s11.data_out;
alias fi_targets[1379] = dv_top.dut.ID.RegFile.registers.s11.we;
alias fi_targets[1380] = dv_top.dut.ID.RegFile.registers.s2.data_in;
alias fi_targets[1381] = dv_top.dut.ID.RegFile.registers.s2.data_out;
alias fi_targets[1382] = dv_top.dut.ID.RegFile.registers.s2.we;
alias fi_targets[1383] = dv_top.dut.ID.RegFile.registers.s3.data_in;
alias fi_targets[1384] = dv_top.dut.ID.RegFile.registers.s3.data_out;
alias fi_targets[1385] = dv_top.dut.ID.RegFile.registers.s3.we;
alias fi_targets[1386] = dv_top.dut.ID.RegFile.registers.s4.data_in;
alias fi_targets[1387] = dv_top.dut.ID.RegFile.registers.s4.data_out;
alias fi_targets[1388] = dv_top.dut.ID.RegFile.registers.s4.we;
alias fi_targets[1389] = dv_top.dut.ID.RegFile.registers.s5.data_in;
alias fi_targets[1390] = dv_top.dut.ID.RegFile.registers.s5.data_out;
alias fi_targets[1391] = dv_top.dut.ID.RegFile.registers.s5.we;
alias fi_targets[1392] = dv_top.dut.ID.RegFile.registers.s6.data_in;
alias fi_targets[1393] = dv_top.dut.ID.RegFile.registers.s6.data_out;
alias fi_targets[1394] = dv_top.dut.ID.RegFile.registers.s6.we;
alias fi_targets[1395] = dv_top.dut.ID.RegFile.registers.s7.data_in;
alias fi_targets[1396] = dv_top.dut.ID.RegFile.registers.s7.data_out;
alias fi_targets[1397] = dv_top.dut.ID.RegFile.registers.s7.we;
alias fi_targets[1398] = dv_top.dut.ID.RegFile.registers.s8.data_in;
alias fi_targets[1399] = dv_top.dut.ID.RegFile.registers.s8.data_out;
alias fi_targets[1400] = dv_top.dut.ID.RegFile.registers.s8.we;
alias fi_targets[1401] = dv_top.dut.ID.RegFile.registers.s9.data_in;
alias fi_targets[1402] = dv_top.dut.ID.RegFile.registers.s9.data_out;
alias fi_targets[1403] = dv_top.dut.ID.RegFile.registers.s9.we;
alias fi_targets[1404] = dv_top.dut.ID.RegFile.registers.sp.data_in;
alias fi_targets[1405] = dv_top.dut.ID.RegFile.registers.sp.data_out;
alias fi_targets[1406] = dv_top.dut.ID.RegFile.registers.sp.we;
alias fi_targets[1407] = dv_top.dut.ID.RegFile.registers.t0.data_in;
alias fi_targets[1408] = dv_top.dut.ID.RegFile.registers.t0.data_out;
alias fi_targets[1409] = dv_top.dut.ID.RegFile.registers.t0.we;
alias fi_targets[1410] = dv_top.dut.ID.RegFile.registers.t1.data_in;
alias fi_targets[1411] = dv_top.dut.ID.RegFile.registers.t1.data_out;
alias fi_targets[1412] = dv_top.dut.ID.RegFile.registers.t1.we;
alias fi_targets[1413] = dv_top.dut.ID.RegFile.registers.t2.data_in;
alias fi_targets[1414] = dv_top.dut.ID.RegFile.registers.t2.data_out;
alias fi_targets[1415] = dv_top.dut.ID.RegFile.registers.t2.we;
alias fi_targets[1416] = dv_top.dut.ID.RegFile.registers.t3.data_in;
alias fi_targets[1417] = dv_top.dut.ID.RegFile.registers.t3.data_out;
alias fi_targets[1418] = dv_top.dut.ID.RegFile.registers.t3.we;
alias fi_targets[1419] = dv_top.dut.ID.RegFile.registers.t4.data_in;
alias fi_targets[1420] = dv_top.dut.ID.RegFile.registers.t4.data_out;
alias fi_targets[1421] = dv_top.dut.ID.RegFile.registers.t4.we;
alias fi_targets[1422] = dv_top.dut.ID.RegFile.registers.t5.data_in;
alias fi_targets[1423] = dv_top.dut.ID.RegFile.registers.t5.data_out;
alias fi_targets[1424] = dv_top.dut.ID.RegFile.registers.t5.we;
alias fi_targets[1425] = dv_top.dut.ID.RegFile.registers.t6.data_in;
alias fi_targets[1426] = dv_top.dut.ID.RegFile.registers.t6.data_out;
alias fi_targets[1427] = dv_top.dut.ID.RegFile.registers.t6.we;
alias fi_targets[1428] = dv_top.dut.ID.RegFile.registers.tp.data_in;
alias fi_targets[1429] = dv_top.dut.ID.RegFile.registers.tp.data_out;
alias fi_targets[1430] = dv_top.dut.ID.RegFile.registers.tp.we;
alias fi_targets[1431] = dv_top.dut.ID.RegFile.registers.zero.data_in;
alias fi_targets[1432] = dv_top.dut.ID.RegFile.registers.zero.data_out;
alias fi_targets[1433] = dv_top.dut.ID.RegFile.registers.zero.we;
alias fi_targets[1434] = dv_top.dut.ID.RegFile.registers.data_in;
alias fi_targets[1435] = dv_top.dut.ID.RegFile.registers.data_out;
alias fi_targets[1436] = dv_top.dut.ID.RegFile.registers.we;
alias fi_targets[1437] = dv_top.dut.ID.RegFile.registers.wr_sel;
alias fi_targets[1438] = dv_top.dut.ID.RegFile.a_out;
alias fi_targets[1439] = dv_top.dut.ID.RegFile.a_select;
alias fi_targets[1440] = dv_top.dut.ID.RegFile.b_out;
alias fi_targets[1441] = dv_top.dut.ID.RegFile.b_select;
alias fi_targets[1442] = dv_top.dut.ID.RegFile.rd_in;
alias fi_targets[1443] = dv_top.dut.ID.RegFile.reg_out;
alias fi_targets[1444] = dv_top.dut.ID.RegFile.we;
alias fi_targets[1445] = dv_top.dut.ID.RegFile.wr_sel;
alias fi_targets[1446] = dv_top.dut.ID.RegFile.write_addr;
alias fi_targets[1447] = dv_top.dut.ID.decoder.a_select;
alias fi_targets[1448] = dv_top.dut.ID.decoder.b_select;
alias fi_targets[1449] = dv_top.dut.ID.decoder.b_type;
alias fi_targets[1450] = dv_top.dut.ID.decoder.branch_sel;
alias fi_targets[1451] = dv_top.dut.ID.decoder.control_word;
alias fi_targets[1452] = dv_top.dut.ID.decoder.d_addr;
alias fi_targets[1453] = dv_top.dut.ID.decoder.func3;
alias fi_targets[1454] = dv_top.dut.ID.decoder.function_select;
alias fi_targets[1455] = dv_top.dut.ID.decoder.i_type;
alias fi_targets[1456] = dv_top.dut.ID.decoder.instruction;
alias fi_targets[1457] = dv_top.dut.ID.decoder.j_type;
alias fi_targets[1458] = dv_top.dut.ID.decoder.jalr;
alias fi_targets[1459] = dv_top.dut.ID.decoder.load;
alias fi_targets[1460] = dv_top.dut.ID.decoder.mem_width_sel;
alias fi_targets[1461] = dv_top.dut.ID.decoder.r_type;
alias fi_targets[1462] = dv_top.dut.ID.decoder.s_type;
alias fi_targets[1463] = dv_top.dut.ID.decoder.save_pc;
alias fi_targets[1464] = dv_top.dut.ID.decoder.u_type;
alias fi_targets[1465] = dv_top.dut.ID.decoder.use_immediate;
alias fi_targets[1466] = dv_top.dut.ID.decoder.we;
alias fi_targets[1467] = dv_top.dut.ID.branch_perediction_i;
alias fi_targets[1468] = dv_top.dut.ID.branch_prediction_internal;
alias fi_targets[1469] = dv_top.dut.ID.branch_prediction_o;
alias fi_targets[1470] = dv_top.dut.ID.branch_sel_internal;
alias fi_targets[1471] = dv_top.dut.ID.branch_sel_o;
alias fi_targets[1472] = dv_top.dut.ID.buble;
alias fi_targets[1473] = dv_top.dut.ID.control_signal_internal;
alias fi_targets[1474] = dv_top.dut.ID.control_signal_o;
alias fi_targets[1475] = dv_top.dut.ID.control_signal_wb;
alias fi_targets[1476] = dv_top.dut.ID.data_a_internal;
alias fi_targets[1477] = dv_top.dut.ID.data_a_o;
alias fi_targets[1478] = dv_top.dut.ID.data_b_internal;
alias fi_targets[1479] = dv_top.dut.ID.data_b_o;
alias fi_targets[1480] = dv_top.dut.ID.data_in_wb;
alias fi_targets[1481] = dv_top.dut.ID.flush;
alias fi_targets[1482] = dv_top.dut.ID.i_instruction;
alias fi_targets[1483] = dv_top.dut.ID.immediate_i;
alias fi_targets[1484] = dv_top.dut.ID.pc_plus_i;
alias fi_targets[1485] = dv_top.dut.ID.pc_plus_internal;
alias fi_targets[1486] = dv_top.dut.ID.pc_plus_o;
alias fi_targets[1487] = dv_top.dut.ID.reg_b_value;
alias fi_targets[1488] = dv_top.dut.ID.rs1_addr;
alias fi_targets[1489] = dv_top.dut.ID.rs2_addr;
alias fi_targets[1490] = dv_top.dut.ID.store_data_internal;
alias fi_targets[1491] = dv_top.dut.ID.store_data_o;
alias fi_targets[1492] = dv_top.dut.Ins_Fetch.PC.correction_mux.addr;
alias fi_targets[1493] = dv_top.dut.Ins_Fetch.PC.correction_mux.data_in;
alias fi_targets[1494] = dv_top.dut.Ins_Fetch.PC.correction_mux.data_out;
alias fi_targets[1495] = dv_top.dut.Ins_Fetch.PC.correction_mux.inner_data;
alias fi_targets[1496] = dv_top.dut.Ins_Fetch.PC.immeadiate_mux.addr;
alias fi_targets[1497] = dv_top.dut.Ins_Fetch.PC.immeadiate_mux.data_in;
alias fi_targets[1498] = dv_top.dut.Ins_Fetch.PC.immeadiate_mux.data_out;
alias fi_targets[1499] = dv_top.dut.Ins_Fetch.PC.immeadiate_mux.inner_data;
alias fi_targets[1500] = dv_top.dut.Ins_Fetch.PC.out_mux.addr;
alias fi_targets[1501] = dv_top.dut.Ins_Fetch.PC.out_mux.data_in;
alias fi_targets[1502] = dv_top.dut.Ins_Fetch.PC.out_mux.data_out;
alias fi_targets[1503] = dv_top.dut.Ins_Fetch.PC.out_mux.inner_data;
alias fi_targets[1504] = dv_top.dut.Ins_Fetch.PC.buble;
alias fi_targets[1505] = dv_top.dut.Ins_Fetch.PC.correct_pc;
alias fi_targets[1506] = dv_top.dut.Ins_Fetch.PC.current_pc;
alias fi_targets[1507] = dv_top.dut.Ins_Fetch.PC.imm_i;
alias fi_targets[1508] = dv_top.dut.Ins_Fetch.PC.inst_addr;
alias fi_targets[1509] = dv_top.dut.Ins_Fetch.PC.instruction_valid;
alias fi_targets[1510] = dv_top.dut.Ins_Fetch.PC.jalr;
alias fi_targets[1511] = dv_top.dut.Ins_Fetch.PC.jump;
alias fi_targets[1512] = dv_top.dut.Ins_Fetch.PC.misprediction;
alias fi_targets[1513] = dv_top.dut.Ins_Fetch.PC.pc_current_val;
alias fi_targets[1514] = dv_top.dut.Ins_Fetch.PC.pc_new_val;
alias fi_targets[1515] = dv_top.dut.Ins_Fetch.PC.pc_plus;
alias fi_targets[1516] = dv_top.dut.Ins_Fetch.PC.pc_plus_four;
alias fi_targets[1517] = dv_top.dut.Ins_Fetch.PC.pc_plus_imm;
alias fi_targets[1518] = dv_top.dut.Ins_Fetch.PC.pc_save;
alias fi_targets[1519] = dv_top.dut.Ins_Fetch.PC.rs1_plus_imm_prediction;
alias fi_targets[1520] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.MUX.addr;
alias fi_targets[1521] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.MUX.data_in;
alias fi_targets[1522] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.MUX.data_out;
alias fi_targets[1523] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.MUX.inner_data;
alias fi_targets[1524] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.b;
alias fi_targets[1525] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.b_imm;
alias fi_targets[1526] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.i_imm;
alias fi_targets[1527] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.imm_o;
alias fi_targets[1528] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.imm_sel;
alias fi_targets[1529] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.instruction;
alias fi_targets[1530] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.j;
alias fi_targets[1531] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.j_imm;
alias fi_targets[1532] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.s;
alias fi_targets[1533] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.s_imm;
alias fi_targets[1534] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.u;
alias fi_targets[1535] = dv_top.dut.Ins_Fetch.early_stage_imm_dec.u_imm;
alias fi_targets[1536] = dv_top.dut.Ins_Fetch.jump_controller.b_type;
alias fi_targets[1537] = dv_top.dut.Ins_Fetch.jump_controller.instruction;
alias fi_targets[1538] = dv_top.dut.Ins_Fetch.jump_controller.j_type;
alias fi_targets[1539] = dv_top.dut.Ins_Fetch.jump_controller.jalr;
alias fi_targets[1540] = dv_top.dut.Ins_Fetch.jump_controller.jump;
alias fi_targets[1541] = dv_top.dut.Ins_Fetch.branch_prediction_o;
alias fi_targets[1542] = dv_top.dut.Ins_Fetch.buble;
alias fi_targets[1543] = dv_top.dut.Ins_Fetch.correct_pc;
alias fi_targets[1544] = dv_top.dut.Ins_Fetch.current_pc;
alias fi_targets[1545] = dv_top.dut.Ins_Fetch.flush;
alias fi_targets[1546] = dv_top.dut.Ins_Fetch.imm;
alias fi_targets[1547] = dv_top.dut.Ins_Fetch.imm_o;
alias fi_targets[1548] = dv_top.dut.Ins_Fetch.inst_addr;
alias fi_targets[1549] = dv_top.dut.Ins_Fetch.instruction_i;
alias fi_targets[1550] = dv_top.dut.Ins_Fetch.instruction_o;
alias fi_targets[1551] = dv_top.dut.Ins_Fetch.instruction_valid;
alias fi_targets[1552] = dv_top.dut.Ins_Fetch.jalr;
alias fi_targets[1553] = dv_top.dut.Ins_Fetch.jump;
alias fi_targets[1554] = dv_top.dut.Ins_Fetch.misprediction;
alias fi_targets[1555] = dv_top.dut.Ins_Fetch.pc_plus_internal;
alias fi_targets[1556] = dv_top.dut.Ins_Fetch.pc_plus_o;
alias fi_targets[1557] = dv_top.dut.MEM.store_data_organizer.MUX_mask1.addr;
alias fi_targets[1558] = dv_top.dut.MEM.store_data_organizer.MUX_mask1.data_in;
alias fi_targets[1559] = dv_top.dut.MEM.store_data_organizer.MUX_mask1.data_out;
alias fi_targets[1560] = dv_top.dut.MEM.store_data_organizer.MUX_mask1.inner_data;
alias fi_targets[1561] = dv_top.dut.MEM.store_data_organizer.MUX_mask2.addr;
alias fi_targets[1562] = dv_top.dut.MEM.store_data_organizer.MUX_mask2.data_in;
alias fi_targets[1563] = dv_top.dut.MEM.store_data_organizer.MUX_mask2.data_out;
alias fi_targets[1564] = dv_top.dut.MEM.store_data_organizer.MUX_mask2.inner_data;
alias fi_targets[1565] = dv_top.dut.MEM.store_data_organizer.Type_sel;
alias fi_targets[1566] = dv_top.dut.MEM.store_data_organizer.data_in;
alias fi_targets[1567] = dv_top.dut.MEM.store_data_organizer.data_out;
alias fi_targets[1568] = dv_top.dut.MEM.store_data_organizer.mask1;
alias fi_targets[1569] = dv_top.dut.MEM.store_data_organizer.mask2;
alias fi_targets[1570] = dv_top.dut.MEM.store_data_organizer.sign;
alias fi_targets[1571] = dv_top.dut.MEM.store_data_organizer.size_sel;
alias fi_targets[1572] = dv_top.dut.MEM.control_signal_i;
alias fi_targets[1573] = dv_top.dut.MEM.control_signal_internal;
alias fi_targets[1574] = dv_top.dut.MEM.control_signal_o;
alias fi_targets[1575] = dv_top.dut.MEM.data_mem_rw;
alias fi_targets[1576] = dv_top.dut.MEM.data_mem_width_sel;
alias fi_targets[1577] = dv_top.dut.MEM.execute_result_i;
alias fi_targets[1578] = dv_top.dut.MEM.execute_result_internal;
alias fi_targets[1579] = dv_top.dut.MEM.execute_result_o;
alias fi_targets[1580] = dv_top.dut.MEM.mem_stage_destination;
alias fi_targets[1581] = dv_top.dut.MEM.mem_stage_we;
alias fi_targets[1582] = dv_top.dut.MEM.store_data_i;
alias fi_targets[1583] = dv_top.dut.MEM.store_data_o;
alias fi_targets[1584] = dv_top.dut.WB.Final_mux.addr;
alias fi_targets[1585] = dv_top.dut.WB.Final_mux.data_in;
alias fi_targets[1586] = dv_top.dut.WB.Final_mux.data_out;
alias fi_targets[1587] = dv_top.dut.WB.Final_mux.inner_data;
alias fi_targets[1588] = dv_top.dut.WB.load_data_organizer.MUX_mask1.addr;
alias fi_targets[1589] = dv_top.dut.WB.load_data_organizer.MUX_mask1.data_in;
alias fi_targets[1590] = dv_top.dut.WB.load_data_organizer.MUX_mask1.data_out;
alias fi_targets[1591] = dv_top.dut.WB.load_data_organizer.MUX_mask1.inner_data;
alias fi_targets[1592] = dv_top.dut.WB.load_data_organizer.MUX_mask2.addr;
alias fi_targets[1593] = dv_top.dut.WB.load_data_organizer.MUX_mask2.data_in;
alias fi_targets[1594] = dv_top.dut.WB.load_data_organizer.MUX_mask2.data_out;
alias fi_targets[1595] = dv_top.dut.WB.load_data_organizer.MUX_mask2.inner_data;
alias fi_targets[1596] = dv_top.dut.WB.load_data_organizer.Type_sel;
alias fi_targets[1597] = dv_top.dut.WB.load_data_organizer.data_in;
alias fi_targets[1598] = dv_top.dut.WB.load_data_organizer.data_out;
alias fi_targets[1599] = dv_top.dut.WB.load_data_organizer.mask1;
alias fi_targets[1600] = dv_top.dut.WB.load_data_organizer.mask2;
alias fi_targets[1601] = dv_top.dut.WB.load_data_organizer.sign;
alias fi_targets[1602] = dv_top.dut.WB.load_data_organizer.size_sel;
alias fi_targets[1603] = dv_top.dut.WB.control_signal_i;
alias fi_targets[1604] = dv_top.dut.WB.control_signal_o;
alias fi_targets[1605] = dv_top.dut.WB.ex_stage_result_i;
alias fi_targets[1606] = dv_top.dut.WB.load_data_i;
alias fi_targets[1607] = dv_top.dut.WB.load_data_internal;
alias fi_targets[1608] = dv_top.dut.WB.wb_result_o;
alias fi_targets[1609] = dv_top.dut.WB.wb_stage_destination;
alias fi_targets[1610] = dv_top.dut.WB.wb_stage_we;
alias fi_targets[1611] = dv_top.dut.A_EX_i;
alias fi_targets[1612] = dv_top.dut.A_sel_DF;
alias fi_targets[1613] = dv_top.dut.B_EX_i;
alias fi_targets[1614] = dv_top.dut.B_sel_DF;
alias fi_targets[1615] = dv_top.dut.Branch_sel_EX_i;
alias fi_targets[1616] = dv_top.dut.Control_Signal_EX_i;
alias fi_targets[1617] = dv_top.dut.Control_Signal_MEM_i;
alias fi_targets[1618] = dv_top.dut.Control_Signal_WB_i;
alias fi_targets[1619] = dv_top.dut.Control_Signal_WB_o;
alias fi_targets[1620] = dv_top.dut.FU_MEM_i;
alias fi_targets[1621] = dv_top.dut.FU_WB_i;
alias fi_targets[1622] = dv_top.dut.Final_Result_WB_o;
alias fi_targets[1623] = dv_top.dut.IMM_ID_i;
alias fi_targets[1624] = dv_top.dut.MEM_result_WB_i;
alias fi_targets[1625] = dv_top.dut.PCPlus_ID_i;
alias fi_targets[1626] = dv_top.dut.PCplus_EX_i;
alias fi_targets[1627] = dv_top.dut.Predicted_MPC_EX_i;
alias fi_targets[1628] = dv_top.dut.Predicted_MPC_ID_i;
alias fi_targets[1629] = dv_top.dut.RAM_DATA_EX_i;
alias fi_targets[1630] = dv_top.dut.RAM_DATA_MEM_i;
alias fi_targets[1631] = dv_top.dut.RA_DF;
alias fi_targets[1632] = dv_top.dut.RB_DF;
alias fi_targets[1633] = dv_top.dut.RD_MEM;
alias fi_targets[1634] = dv_top.dut.RD_WB;
alias fi_targets[1635] = dv_top.dut.WE_MEM;
alias fi_targets[1636] = dv_top.dut.WE_WB;
alias fi_targets[1637] = dv_top.dut.buble;
alias fi_targets[1638] = dv_top.dut.correct_pc;
alias fi_targets[1639] = dv_top.dut.data_mem_addr_o;
alias fi_targets[1640] = dv_top.dut.data_mem_control;
alias fi_targets[1641] = dv_top.dut.data_mem_data_rd_data;
alias fi_targets[1642] = dv_top.dut.data_mem_data_wr_data;
alias fi_targets[1643] = dv_top.dut.data_mem_rw;
alias fi_targets[1644] = dv_top.dut.ins_address;
alias fi_targets[1645] = dv_top.dut.instruction_ID_i;
alias fi_targets[1646] = dv_top.dut.instruction_i;
alias fi_targets[1647] = dv_top.dut.instruction_valid;
alias fi_targets[1648] = dv_top.dut.misprediction;
alias fi_targets[1649] = dv_top.dut.rs1_id;
alias fi_targets[1650] = dv_top.dut.rs2_id;
alias fi_targets[1651] = dv_top.dut.store_sel_df;